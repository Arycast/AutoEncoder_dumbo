library verilog;
use verilog.vl_types.all;
entity top_level_architecture is
    port(
        clock           : in     vl_logic
    );
end top_level_architecture;
