library verilog;
use verilog.vl_types.all;
entity ALU_cells is
    port(
        input_mem_1_1   : in     vl_logic_vector(15 downto 0);
        input_mem_1_2   : in     vl_logic_vector(15 downto 0);
        input_mem_1_3   : in     vl_logic_vector(15 downto 0);
        input_mem_1_4   : in     vl_logic_vector(15 downto 0);
        input_mem_1_5   : in     vl_logic_vector(15 downto 0);
        input_mem_1_6   : in     vl_logic_vector(15 downto 0);
        input_mem_1_7   : in     vl_logic_vector(15 downto 0);
        input_mem_1_8   : in     vl_logic_vector(15 downto 0);
        input_mem_1_9   : in     vl_logic_vector(15 downto 0);
        input_mem_2_1   : in     vl_logic_vector(15 downto 0);
        input_mem_2_2   : in     vl_logic_vector(15 downto 0);
        input_mem_2_3   : in     vl_logic_vector(15 downto 0);
        input_mem_2_4   : in     vl_logic_vector(15 downto 0);
        input_mem_2_5   : in     vl_logic_vector(15 downto 0);
        input_mem_2_6   : in     vl_logic_vector(15 downto 0);
        input_mem_2_7   : in     vl_logic_vector(15 downto 0);
        input_mem_2_8   : in     vl_logic_vector(15 downto 0);
        input_mem_2_9   : in     vl_logic_vector(15 downto 0);
        input_weight    : in     vl_logic_vector(15 downto 0);
        input_bias      : in     vl_logic_vector(15 downto 0);
        output_bias     : in     vl_logic_vector(15 downto 0);
        output_error    : in     vl_logic_vector(15 downto 0);
        output_weight_diff: in     vl_logic_vector(15 downto 0);
        input_weight_diff: in     vl_logic_vector(15 downto 0);
        middle_layer_error: in     vl_logic_vector(15 downto 0);
        output_pixel    : in     vl_logic_vector(15 downto 0);
        input_pixel     : in     vl_logic_vector(15 downto 0);
        mux_1_control   : in     vl_logic_vector(4 downto 0);
        mux_2_control   : in     vl_logic_vector(4 downto 0);
        mux_3_control   : in     vl_logic_vector(1 downto 0);
        mux_4_control   : in     vl_logic_vector(3 downto 0);
        enable_ALU      : in     vl_logic;
        op_select       : in     vl_logic_vector(1 downto 0);
        demux_1_control : in     vl_logic_vector(3 downto 0);
        to_memory       : out    vl_logic_vector(15 downto 0);
        to_sigmoid      : out    vl_logic_vector(15 downto 0);
        to_input_weight : out    vl_logic_vector(15 downto 0);
        to_input_bias   : out    vl_logic_vector(15 downto 0);
        to_output_bias  : out    vl_logic_vector(15 downto 0);
        to_output_error : out    vl_logic_vector(15 downto 0);
        to_output_weight_diff: out    vl_logic_vector(15 downto 0);
        to_input_weight_diff: out    vl_logic_vector(15 downto 0);
        to_middle_layer_error: out    vl_logic_vector(15 downto 0)
    );
end ALU_cells;
