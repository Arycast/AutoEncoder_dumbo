<<<<<<< HEAD
//////////////////////////////////////////////////////////////////////////////////
// Engineer    : Achmad novel, Fauzan Ibrahim, Nicholas Teffandi
// Design Name : Autoencoder
// Module Name : sigmoid_lut
// Project Name: Autoencoder
//////////////////////////////////////////////////////////////////////////////////

// Input and Output is Unsigned

module sigmoid_lut (
   input wire [15:0] addr,
   output reg [15:0] result
);

   always @(*) begin
      
      case (addr)
         63744    :	result = 16'd0;
         63745    :	result = 16'd0;
         63746    :	result = 16'd0;
         63747    :	result = 16'd0;
         63748    :	result = 16'd0;
         63749    :	result = 16'd0;
         63750    :	result = 16'd0;
         63751    :	result = 16'd0;
         63752    :	result = 16'd0;
         63753    :	result = 16'd0;
         63754    :	result = 16'd0;
         63755    :	result = 16'd0;
         63756    :	result = 16'd0;
         63757    :	result = 16'd0;
         63758    :	result = 16'd0;
         63759    :	result = 16'd0;
         63760    :	result = 16'd0;
         63761    :	result = 16'd0;
         63762    :	result = 16'd0;
         63763    :	result = 16'd0;
         63764    :	result = 16'd0;
         63765    :	result = 16'd0;
         63766    :	result = 16'd0;
         63767    :	result = 16'd0;
         63768    :	result = 16'd0;
         63769    :	result = 16'd0;
         63770    :	result = 16'd0;
         63771    :	result = 16'd0;
         63772    :	result = 16'd0;
         63773    :	result = 16'd0;
         63774    :	result = 16'd0;
         63775    :	result = 16'd0;
         63776    :	result = 16'd0;
         63777    :	result = 16'd0;
         63778    :	result = 16'd0;
         63779    :	result = 16'd0;
         63780    :	result = 16'd0;
         63781    :	result = 16'd0;
         63782    :	result = 16'd0;
         63783    :	result = 16'd0;
         63784    :	result = 16'd0;
         63785    :	result = 16'd0;
         63786    :	result = 16'd0;
         63787    :	result = 16'd0;
         63788    :	result = 16'd0;
         63789    :	result = 16'd0;
         63790    :	result = 16'd0;
         63791    :	result = 16'd0;
         63792    :	result = 16'd0;
         63793    :	result = 16'd0;
         63794    :	result = 16'd0;
         63795    :	result = 16'd0;
         63796    :	result = 16'd0;
         63797    :	result = 16'd0;
         63798    :	result = 16'd0;
         63799    :	result = 16'd0;
         63800    :	result = 16'd0;
         63801    :	result = 16'd0;
         63802    :	result = 16'd0;
         63803    :	result = 16'd0;
         63804    :	result = 16'd0;
         63805    :	result = 16'd0;
         63806    :	result = 16'd0;
         63807    :	result = 16'd0;
         63808    :	result = 16'd0;
         63809    :	result = 16'd0;
         63810    :	result = 16'd0;
         63811    :	result = 16'd0;
         63812    :	result = 16'd0;
         63813    :	result = 16'd0;
         63814    :	result = 16'd0;
         63815    :	result = 16'd0;
         63816    :	result = 16'd0;
         63817    :	result = 16'd0;
         63818    :	result = 16'd0;
         63819    :	result = 16'd0;
         63820    :	result = 16'd0;
         63821    :	result = 16'd0;
         63822    :	result = 16'd0;
         63823    :	result = 16'd0;
         63824    :	result = 16'd0;
         63825    :	result = 16'd0;
         63826    :	result = 16'd0;
         63827    :	result = 16'd0;
         63828    :	result = 16'd0;
         63829    :	result = 16'd0;
         63830    :	result = 16'd0;
         63831    :	result = 16'd0;
         63832    :	result = 16'd0;
         63833    :	result = 16'd0;
         63834    :	result = 16'd0;
         63835    :	result = 16'd0;
         63836    :	result = 16'd0;
         63837    :	result = 16'd0;
         63838    :	result = 16'd0;
         63839    :	result = 16'd0;
         63840    :	result = 16'd0;
         63841    :	result = 16'd0;
         63842    :	result = 16'd0;
         63843    :	result = 16'd0;
         63844    :	result = 16'd0;
         63845    :	result = 16'd0;
         63846    :	result = 16'd0;
         63847    :	result = 16'd0;
         63848    :	result = 16'd0;
         63849    :	result = 16'd0;
         63850    :	result = 16'd0;
         63851    :	result = 16'd0;
         63852    :	result = 16'd0;
         63853    :	result = 16'd0;
         63854    :	result = 16'd0;
         63855    :	result = 16'd0;
         63856    :	result = 16'd0;
         63857    :	result = 16'd0;
         63858    :	result = 16'd0;
         63859    :	result = 16'd0;
         63860    :	result = 16'd0;
         63861    :	result = 16'd0;
         63862    :	result = 16'd0;
         63863    :	result = 16'd0;
         63864    :	result = 16'd0;
         63865    :	result = 16'd0;
         63866    :	result = 16'd0;
         63867    :	result = 16'd0;
         63868    :	result = 16'd0;
         63869    :	result = 16'd0;
         63870    :	result = 16'd0;
         63871    :	result = 16'd0;
         63872    :	result = 16'd0;
         63873    :	result = 16'd0;
         63874    :	result = 16'd0;
         63875    :	result = 16'd0;
         63876    :	result = 16'd0;
         63877    :	result = 16'd0;
         63878    :	result = 16'd0;
         63879    :	result = 16'd0;
         63880    :	result = 16'd0;
         63881    :	result = 16'd0;
         63882    :	result = 16'd0;
         63883    :	result = 16'd0;
         63884    :	result = 16'd0;
         63885    :	result = 16'd0;
         63886    :	result = 16'd0;
         63887    :	result = 16'd0;
         63888    :	result = 16'd0;
         63889    :	result = 16'd0;
         63890    :	result = 16'd0;
         63891    :	result = 16'd0;
         63892    :	result = 16'd0;
         63893    :	result = 16'd0;
         63894    :	result = 16'd0;
         63895    :	result = 16'd0;
         63896    :	result = 16'd0;
         63897    :	result = 16'd0;
         63898    :	result = 16'd0;
         63899    :	result = 16'd0;
         63900    :	result = 16'd0;
         63901    :	result = 16'd0;
         63902    :	result = 16'd0;
         63903    :	result = 16'd0;
         63904    :	result = 16'd0;
         63905    :	result = 16'd0;
         63906    :	result = 16'd0;
         63907    :	result = 16'd0;
         63908    :	result = 16'd0;
         63909    :	result = 16'd0;
         63910    :	result = 16'd0;
         63911    :	result = 16'd0;
         63912    :	result = 16'd0;
         63913    :	result = 16'd0;
         63914    :	result = 16'd0;
         63915    :	result = 16'd0;
         63916    :	result = 16'd0;
         63917    :	result = 16'd0;
         63918    :	result = 16'd0;
         63919    :	result = 16'd0;
         63920    :	result = 16'd0;
         63921    :	result = 16'd0;
         63922    :	result = 16'd0;
         63923    :	result = 16'd0;
         63924    :	result = 16'd0;
         63925    :	result = 16'd0;
         63926    :	result = 16'd0;
         63927    :	result = 16'd0;
         63928    :	result = 16'd0;
         63929    :	result = 16'd0;
         63930    :	result = 16'd0;
         63931    :	result = 16'd0;
         63932    :	result = 16'd0;
         63933    :	result = 16'd0;
         63934    :	result = 16'd0;
         63935    :	result = 16'd0;
         63936    :	result = 16'd0;
         63937    :	result = 16'd0;
         63938    :	result = 16'd0;
         63939    :	result = 16'd0;
         63940    :	result = 16'd0;
         63941    :	result = 16'd0;
         63942    :	result = 16'd0;
         63943    :	result = 16'd0;
         63944    :	result = 16'd0;
         63945    :	result = 16'd0;
         63946    :	result = 16'd0;
         63947    :	result = 16'd0;
         63948    :	result = 16'd0;
         63949    :	result = 16'd0;
         63950    :	result = 16'd0;
         63951    :	result = 16'd0;
         63952    :	result = 16'd0;
         63953    :	result = 16'd0;
         63954    :	result = 16'd0;
         63955    :	result = 16'd0;
         63956    :	result = 16'd0;
         63957    :	result = 16'd0;
         63958    :	result = 16'd0;
         63959    :	result = 16'd0;
         63960    :	result = 16'd0;
         63961    :	result = 16'd0;
         63962    :	result = 16'd0;
         63963    :	result = 16'd0;
         63964    :	result = 16'd0;
         63965    :	result = 16'd0;
         63966    :	result = 16'd0;
         63967    :	result = 16'd0;
         63968    :	result = 16'd0;
         63969    :	result = 16'd0;
         63970    :	result = 16'd0;
         63971    :	result = 16'd0;
         63972    :	result = 16'd0;
         63973    :	result = 16'd0;
         63974    :	result = 16'd0;
         63975    :	result = 16'd0;
         63976    :	result = 16'd0;
         63977    :	result = 16'd0;
         63978    :	result = 16'd0;
         63979    :	result = 16'd0;
         63980    :	result = 16'd0;
         63981    :	result = 16'd0;
         63982    :	result = 16'd0;
         63983    :	result = 16'd0;
         63984    :	result = 16'd0;
         63985    :	result = 16'd0;
         63986    :	result = 16'd0;
         63987    :	result = 16'd0;
         63988    :	result = 16'd0;
         63989    :	result = 16'd0;
         63990    :	result = 16'd0;
         63991    :	result = 16'd0;
         63992    :	result = 16'd0;
         63993    :	result = 16'd0;
         63994    :	result = 16'd0;
         63995    :	result = 16'd0;
         63996    :	result = 16'd0;
         63997    :	result = 16'd0;
         63998    :	result = 16'd0;
         63999    :	result = 16'd0;
         64000    :	result = 16'd0;
         64001    :	result = 16'd0;
         64002    :	result = 16'd0;
         64003    :	result = 16'd0;
         64004    :	result = 16'd0;
         64005    :	result = 16'd0;
         64006    :	result = 16'd0;
         64007    :	result = 16'd0;
         64008    :	result = 16'd0;
         64009    :	result = 16'd0;
         64010    :	result = 16'd0;
         64011    :	result = 16'd0;
         64012    :	result = 16'd0;
         64013    :	result = 16'd0;
         64014    :	result = 16'd0;
         64015    :	result = 16'd0;
         64016    :	result = 16'd0;
         64017    :	result = 16'd0;
         64018    :	result = 16'd0;
         64019    :	result = 16'd0;
         64020    :	result = 16'd0;
         64021    :	result = 16'd0;
         64022    :	result = 16'd0;
         64023    :	result = 16'd0;
         64024    :	result = 16'd0;
         64025    :	result = 16'd0;
         64026    :	result = 16'd0;
         64027    :	result = 16'd0;
         64028    :	result = 16'd0;
         64029    :	result = 16'd0;
         64030    :	result = 16'd0;
         64031    :	result = 16'd0;
         64032    :	result = 16'd0;
         64033    :	result = 16'd0;
         64034    :	result = 16'd0;
         64035    :	result = 16'd0;
         64036    :	result = 16'd0;
         64037    :	result = 16'd0;
         64038    :	result = 16'd0;
         64039    :	result = 16'd0;
         64040    :	result = 16'd0;
         64041    :	result = 16'd0;
         64042    :	result = 16'd0;
         64043    :	result = 16'd0;
         64044    :	result = 16'd0;
         64045    :	result = 16'd0;
         64046    :	result = 16'd0;
         64047    :	result = 16'd0;
         64048    :	result = 16'd0;
         64049    :	result = 16'd0;
         64050    :	result = 16'd0;
         64051    :	result = 16'd0;
         64052    :	result = 16'd0;
         64053    :	result = 16'd0;
         64054    :	result = 16'd0;
         64055    :	result = 16'd0;
         64056    :	result = 16'd0;
         64057    :	result = 16'd0;
         64058    :	result = 16'd0;
         64059    :	result = 16'd0;
         64060    :	result = 16'd0;
         64061    :	result = 16'd0;
         64062    :	result = 16'd0;
         64063    :	result = 16'd0;
         64064    :	result = 16'd0;
         64065    :	result = 16'd0;
         64066    :	result = 16'd0;
         64067    :	result = 16'd0;
         64068    :	result = 16'd0;
         64069    :	result = 16'd0;
         64070    :	result = 16'd0;
         64071    :	result = 16'd0;
         64072    :	result = 16'd0;
         64073    :	result = 16'd0;
         64074    :	result = 16'd0;
         64075    :	result = 16'd0;
         64076    :	result = 16'd0;
         64077    :	result = 16'd0;
         64078    :	result = 16'd0;
         64079    :	result = 16'd0;
         64080    :	result = 16'd0;
         64081    :	result = 16'd0;
         64082    :	result = 16'd0;
         64083    :	result = 16'd0;
         64084    :	result = 16'd0;
         64085    :	result = 16'd0;
         64086    :	result = 16'd0;
         64087    :	result = 16'd0;
         64088    :	result = 16'd0;
         64089    :	result = 16'd0;
         64090    :	result = 16'd0;
         64091    :	result = 16'd0;
         64092    :	result = 16'd0;
         64093    :	result = 16'd0;
         64094    :	result = 16'd0;
         64095    :	result = 16'd0;
         64096    :	result = 16'd0;
         64097    :	result = 16'd0;
         64098    :	result = 16'd0;
         64099    :	result = 16'd0;
         64100    :	result = 16'd0;
         64101    :	result = 16'd0;
         64102    :	result = 16'd0;
         64103    :	result = 16'd0;
         64104    :	result = 16'd0;
         64105    :	result = 16'd0;
         64106    :	result = 16'd0;
         64107    :	result = 16'd0;
         64108    :	result = 16'd0;
         64109    :	result = 16'd0;
         64110    :	result = 16'd0;
         64111    :	result = 16'd0;
         64112    :	result = 16'd0;
         64113    :	result = 16'd0;
         64114    :	result = 16'd0;
         64115    :	result = 16'd0;
         64116    :	result = 16'd0;
         64117    :	result = 16'd1;
         64118    :	result = 16'd1;
         64119    :	result = 16'd1;
         64120    :	result = 16'd1;
         64121    :	result = 16'd1;
         64122    :	result = 16'd1;
         64123    :	result = 16'd1;
         64124    :	result = 16'd1;
         64125    :	result = 16'd1;
         64126    :	result = 16'd1;
         64127    :	result = 16'd1;
         64128    :	result = 16'd1;
         64129    :	result = 16'd1;
         64130    :	result = 16'd1;
         64131    :	result = 16'd1;
         64132    :	result = 16'd1;
         64133    :	result = 16'd1;
         64134    :	result = 16'd1;
         64135    :	result = 16'd1;
         64136    :	result = 16'd1;
         64137    :	result = 16'd1;
         64138    :	result = 16'd1;
         64139    :	result = 16'd1;
         64140    :	result = 16'd1;
         64141    :	result = 16'd1;
         64142    :	result = 16'd1;
         64143    :	result = 16'd1;
         64144    :	result = 16'd1;
         64145    :	result = 16'd1;
         64146    :	result = 16'd1;
         64147    :	result = 16'd1;
         64148    :	result = 16'd1;
         64149    :	result = 16'd1;
         64150    :	result = 16'd1;
         64151    :	result = 16'd1;
         64152    :	result = 16'd1;
         64153    :	result = 16'd1;
         64154    :	result = 16'd1;
         64155    :	result = 16'd1;
         64156    :	result = 16'd1;
         64157    :	result = 16'd1;
         64158    :	result = 16'd1;
         64159    :	result = 16'd1;
         64160    :	result = 16'd1;
         64161    :	result = 16'd1;
         64162    :	result = 16'd1;
         64163    :	result = 16'd1;
         64164    :	result = 16'd1;
         64165    :	result = 16'd1;
         64166    :	result = 16'd1;
         64167    :	result = 16'd1;
         64168    :	result = 16'd1;
         64169    :	result = 16'd1;
         64170    :	result = 16'd1;
         64171    :	result = 16'd1;
         64172    :	result = 16'd1;
         64173    :	result = 16'd1;
         64174    :	result = 16'd1;
         64175    :	result = 16'd1;
         64176    :	result = 16'd1;
         64177    :	result = 16'd1;
         64178    :	result = 16'd1;
         64179    :	result = 16'd1;
         64180    :	result = 16'd1;
         64181    :	result = 16'd1;
         64182    :	result = 16'd1;
         64183    :	result = 16'd1;
         64184    :	result = 16'd1;
         64185    :	result = 16'd1;
         64186    :	result = 16'd1;
         64187    :	result = 16'd1;
         64188    :	result = 16'd1;
         64189    :	result = 16'd1;
         64190    :	result = 16'd1;
         64191    :	result = 16'd1;
         64192    :	result = 16'd1;
         64193    :	result = 16'd1;
         64194    :	result = 16'd1;
         64195    :	result = 16'd1;
         64196    :	result = 16'd1;
         64197    :	result = 16'd1;
         64198    :	result = 16'd1;
         64199    :	result = 16'd1;
         64200    :	result = 16'd1;
         64201    :	result = 16'd1;
         64202    :	result = 16'd1;
         64203    :	result = 16'd1;
         64204    :	result = 16'd1;
         64205    :	result = 16'd1;
         64206    :	result = 16'd1;
         64207    :	result = 16'd1;
         64208    :	result = 16'd1;
         64209    :	result = 16'd1;
         64210    :	result = 16'd1;
         64211    :	result = 16'd1;
         64212    :	result = 16'd1;
         64213    :	result = 16'd1;
         64214    :	result = 16'd1;
         64215    :	result = 16'd1;
         64216    :	result = 16'd1;
         64217    :	result = 16'd1;
         64218    :	result = 16'd1;
         64219    :	result = 16'd1;
         64220    :	result = 16'd1;
         64221    :	result = 16'd1;
         64222    :	result = 16'd1;
         64223    :	result = 16'd1;
         64224    :	result = 16'd1;
         64225    :	result = 16'd1;
         64226    :	result = 16'd1;
         64227    :	result = 16'd1;
         64228    :	result = 16'd1;
         64229    :	result = 16'd1;
         64230    :	result = 16'd1;
         64231    :	result = 16'd1;
         64232    :	result = 16'd1;
         64233    :	result = 16'd1;
         64234    :	result = 16'd1;
         64235    :	result = 16'd1;
         64236    :	result = 16'd1;
         64237    :	result = 16'd1;
         64238    :	result = 16'd1;
         64239    :	result = 16'd1;
         64240    :	result = 16'd1;
         64241    :	result = 16'd1;
         64242    :	result = 16'd1;
         64243    :	result = 16'd1;
         64244    :	result = 16'd1;
         64245    :	result = 16'd1;
         64246    :	result = 16'd1;
         64247    :	result = 16'd1;
         64248    :	result = 16'd1;
         64249    :	result = 16'd1;
         64250    :	result = 16'd1;
         64251    :	result = 16'd1;
         64252    :	result = 16'd1;
         64253    :	result = 16'd1;
         64254    :	result = 16'd1;
         64255    :	result = 16'd1;
         64256    :	result = 16'd1;
         64257    :	result = 16'd1;
         64258    :	result = 16'd1;
         64259    :	result = 16'd1;
         64260    :	result = 16'd1;
         64261    :	result = 16'd1;
         64262    :	result = 16'd1;
         64263    :	result = 16'd1;
         64264    :	result = 16'd1;
         64265    :	result = 16'd1;
         64266    :	result = 16'd1;
         64267    :	result = 16'd1;
         64268    :	result = 16'd1;
         64269    :	result = 16'd1;
         64270    :	result = 16'd1;
         64271    :	result = 16'd1;
         64272    :	result = 16'd1;
         64273    :	result = 16'd1;
         64274    :	result = 16'd1;
         64275    :	result = 16'd1;
         64276    :	result = 16'd1;
         64277    :	result = 16'd1;
         64278    :	result = 16'd1;
         64279    :	result = 16'd1;
         64280    :	result = 16'd1;
         64281    :	result = 16'd1;
         64282    :	result = 16'd1;
         64283    :	result = 16'd1;
         64284    :	result = 16'd1;
         64285    :	result = 16'd1;
         64286    :	result = 16'd1;
         64287    :	result = 16'd1;
         64288    :	result = 16'd1;
         64289    :	result = 16'd1;
         64290    :	result = 16'd1;
         64291    :	result = 16'd1;
         64292    :	result = 16'd1;
         64293    :	result = 16'd1;
         64294    :	result = 16'd1;
         64295    :	result = 16'd2;
         64296    :	result = 16'd2;
         64297    :	result = 16'd2;
         64298    :	result = 16'd2;
         64299    :	result = 16'd2;
         64300    :	result = 16'd2;
         64301    :	result = 16'd2;
         64302    :	result = 16'd2;
         64303    :	result = 16'd2;
         64304    :	result = 16'd2;
         64305    :	result = 16'd2;
         64306    :	result = 16'd2;
         64307    :	result = 16'd2;
         64308    :	result = 16'd2;
         64309    :	result = 16'd2;
         64310    :	result = 16'd2;
         64311    :	result = 16'd2;
         64312    :	result = 16'd2;
         64313    :	result = 16'd2;
         64314    :	result = 16'd2;
         64315    :	result = 16'd2;
         64316    :	result = 16'd2;
         64317    :	result = 16'd2;
         64318    :	result = 16'd2;
         64319    :	result = 16'd2;
         64320    :	result = 16'd2;
         64321    :	result = 16'd2;
         64322    :	result = 16'd2;
         64323    :	result = 16'd2;
         64324    :	result = 16'd2;
         64325    :	result = 16'd2;
         64326    :	result = 16'd2;
         64327    :	result = 16'd2;
         64328    :	result = 16'd2;
         64329    :	result = 16'd2;
         64330    :	result = 16'd2;
         64331    :	result = 16'd2;
         64332    :	result = 16'd2;
         64333    :	result = 16'd2;
         64334    :	result = 16'd2;
         64335    :	result = 16'd2;
         64336    :	result = 16'd2;
         64337    :	result = 16'd2;
         64338    :	result = 16'd2;
         64339    :	result = 16'd2;
         64340    :	result = 16'd2;
         64341    :	result = 16'd2;
         64342    :	result = 16'd2;
         64343    :	result = 16'd2;
         64344    :	result = 16'd2;
         64345    :	result = 16'd2;
         64346    :	result = 16'd2;
         64347    :	result = 16'd2;
         64348    :	result = 16'd2;
         64349    :	result = 16'd2;
         64350    :	result = 16'd2;
         64351    :	result = 16'd2;
         64352    :	result = 16'd2;
         64353    :	result = 16'd2;
         64354    :	result = 16'd2;
         64355    :	result = 16'd2;
         64356    :	result = 16'd2;
         64357    :	result = 16'd2;
         64358    :	result = 16'd2;
         64359    :	result = 16'd2;
         64360    :	result = 16'd2;
         64361    :	result = 16'd2;
         64362    :	result = 16'd2;
         64363    :	result = 16'd2;
         64364    :	result = 16'd2;
         64365    :	result = 16'd2;
         64366    :	result = 16'd2;
         64367    :	result = 16'd2;
         64368    :	result = 16'd2;
         64369    :	result = 16'd2;
         64370    :	result = 16'd2;
         64371    :	result = 16'd2;
         64372    :	result = 16'd2;
         64373    :	result = 16'd2;
         64374    :	result = 16'd2;
         64375    :	result = 16'd2;
         64376    :	result = 16'd2;
         64377    :	result = 16'd2;
         64378    :	result = 16'd2;
         64379    :	result = 16'd2;
         64380    :	result = 16'd2;
         64381    :	result = 16'd2;
         64382    :	result = 16'd2;
         64383    :	result = 16'd2;
         64384    :	result = 16'd2;
         64385    :	result = 16'd2;
         64386    :	result = 16'd2;
         64387    :	result = 16'd2;
         64388    :	result = 16'd2;
         64389    :	result = 16'd2;
         64390    :	result = 16'd2;
         64391    :	result = 16'd2;
         64392    :	result = 16'd2;
         64393    :	result = 16'd2;
         64394    :	result = 16'd2;
         64395    :	result = 16'd2;
         64396    :	result = 16'd2;
         64397    :	result = 16'd2;
         64398    :	result = 16'd2;
         64399    :	result = 16'd2;
         64400    :	result = 16'd3;
         64401    :	result = 16'd3;
         64402    :	result = 16'd3;
         64403    :	result = 16'd3;
         64404    :	result = 16'd3;
         64405    :	result = 16'd3;
         64406    :	result = 16'd3;
         64407    :	result = 16'd3;
         64408    :	result = 16'd3;
         64409    :	result = 16'd3;
         64410    :	result = 16'd3;
         64411    :	result = 16'd3;
         64412    :	result = 16'd3;
         64413    :	result = 16'd3;
         64414    :	result = 16'd3;
         64415    :	result = 16'd3;
         64416    :	result = 16'd3;
         64417    :	result = 16'd3;
         64418    :	result = 16'd3;
         64419    :	result = 16'd3;
         64420    :	result = 16'd3;
         64421    :	result = 16'd3;
         64422    :	result = 16'd3;
         64423    :	result = 16'd3;
         64424    :	result = 16'd3;
         64425    :	result = 16'd3;
         64426    :	result = 16'd3;
         64427    :	result = 16'd3;
         64428    :	result = 16'd3;
         64429    :	result = 16'd3;
         64430    :	result = 16'd3;
         64431    :	result = 16'd3;
         64432    :	result = 16'd3;
         64433    :	result = 16'd3;
         64434    :	result = 16'd3;
         64435    :	result = 16'd3;
         64436    :	result = 16'd3;
         64437    :	result = 16'd3;
         64438    :	result = 16'd3;
         64439    :	result = 16'd3;
         64440    :	result = 16'd3;
         64441    :	result = 16'd3;
         64442    :	result = 16'd3;
         64443    :	result = 16'd3;
         64444    :	result = 16'd3;
         64445    :	result = 16'd3;
         64446    :	result = 16'd3;
         64447    :	result = 16'd3;
         64448    :	result = 16'd3;
         64449    :	result = 16'd3;
         64450    :	result = 16'd3;
         64451    :	result = 16'd3;
         64452    :	result = 16'd3;
         64453    :	result = 16'd3;
         64454    :	result = 16'd3;
         64455    :	result = 16'd3;
         64456    :	result = 16'd3;
         64457    :	result = 16'd3;
         64458    :	result = 16'd3;
         64459    :	result = 16'd3;
         64460    :	result = 16'd3;
         64461    :	result = 16'd3;
         64462    :	result = 16'd3;
         64463    :	result = 16'd3;
         64464    :	result = 16'd3;
         64465    :	result = 16'd3;
         64466    :	result = 16'd3;
         64467    :	result = 16'd3;
         64468    :	result = 16'd3;
         64469    :	result = 16'd3;
         64470    :	result = 16'd3;
         64471    :	result = 16'd3;
         64472    :	result = 16'd3;
         64473    :	result = 16'd3;
         64474    :	result = 16'd3;
         64475    :	result = 16'd4;
         64476    :	result = 16'd4;
         64477    :	result = 16'd4;
         64478    :	result = 16'd4;
         64479    :	result = 16'd4;
         64480    :	result = 16'd4;
         64481    :	result = 16'd4;
         64482    :	result = 16'd4;
         64483    :	result = 16'd4;
         64484    :	result = 16'd4;
         64485    :	result = 16'd4;
         64486    :	result = 16'd4;
         64487    :	result = 16'd4;
         64488    :	result = 16'd4;
         64489    :	result = 16'd4;
         64490    :	result = 16'd4;
         64491    :	result = 16'd4;
         64492    :	result = 16'd4;
         64493    :	result = 16'd4;
         64494    :	result = 16'd4;
         64495    :	result = 16'd4;
         64496    :	result = 16'd4;
         64497    :	result = 16'd4;
         64498    :	result = 16'd4;
         64499    :	result = 16'd4;
         64500    :	result = 16'd4;
         64501    :	result = 16'd4;
         64502    :	result = 16'd4;
         64503    :	result = 16'd4;
         64504    :	result = 16'd4;
         64505    :	result = 16'd4;
         64506    :	result = 16'd4;
         64507    :	result = 16'd4;
         64508    :	result = 16'd4;
         64509    :	result = 16'd4;
         64510    :	result = 16'd4;
         64511    :	result = 16'd4;
         64512    :	result = 16'd4;
         64513    :	result = 16'd4;
         64514    :	result = 16'd4;
         64515    :	result = 16'd4;
         64516    :	result = 16'd4;
         64517    :	result = 16'd4;
         64518    :	result = 16'd4;
         64519    :	result = 16'd4;
         64520    :	result = 16'd4;
         64521    :	result = 16'd4;
         64522    :	result = 16'd4;
         64523    :	result = 16'd4;
         64524    :	result = 16'd4;
         64525    :	result = 16'd4;
         64526    :	result = 16'd4;
         64527    :	result = 16'd4;
         64528    :	result = 16'd4;
         64529    :	result = 16'd4;
         64530    :	result = 16'd4;
         64531    :	result = 16'd4;
         64532    :	result = 16'd4;
         64533    :	result = 16'd5;
         64534    :	result = 16'd5;
         64535    :	result = 16'd5;
         64536    :	result = 16'd5;
         64537    :	result = 16'd5;
         64538    :	result = 16'd5;
         64539    :	result = 16'd5;
         64540    :	result = 16'd5;
         64541    :	result = 16'd5;
         64542    :	result = 16'd5;
         64543    :	result = 16'd5;
         64544    :	result = 16'd5;
         64545    :	result = 16'd5;
         64546    :	result = 16'd5;
         64547    :	result = 16'd5;
         64548    :	result = 16'd5;
         64549    :	result = 16'd5;
         64550    :	result = 16'd5;
         64551    :	result = 16'd5;
         64552    :	result = 16'd5;
         64553    :	result = 16'd5;
         64554    :	result = 16'd5;
         64555    :	result = 16'd5;
         64556    :	result = 16'd5;
         64557    :	result = 16'd5;
         64558    :	result = 16'd5;
         64559    :	result = 16'd5;
         64560    :	result = 16'd5;
         64561    :	result = 16'd5;
         64562    :	result = 16'd5;
         64563    :	result = 16'd5;
         64564    :	result = 16'd5;
         64565    :	result = 16'd5;
         64566    :	result = 16'd5;
         64567    :	result = 16'd5;
         64568    :	result = 16'd5;
         64569    :	result = 16'd5;
         64570    :	result = 16'd5;
         64571    :	result = 16'd5;
         64572    :	result = 16'd5;
         64573    :	result = 16'd5;
         64574    :	result = 16'd5;
         64575    :	result = 16'd5;
         64576    :	result = 16'd5;
         64577    :	result = 16'd5;
         64578    :	result = 16'd5;
         64579    :	result = 16'd5;
         64580    :	result = 16'd5;
         64581    :	result = 16'd6;
         64582    :	result = 16'd6;
         64583    :	result = 16'd6;
         64584    :	result = 16'd6;
         64585    :	result = 16'd6;
         64586    :	result = 16'd6;
         64587    :	result = 16'd6;
         64588    :	result = 16'd6;
         64589    :	result = 16'd6;
         64590    :	result = 16'd6;
         64591    :	result = 16'd6;
         64592    :	result = 16'd6;
         64593    :	result = 16'd6;
         64594    :	result = 16'd6;
         64595    :	result = 16'd6;
         64596    :	result = 16'd6;
         64597    :	result = 16'd6;
         64598    :	result = 16'd6;
         64599    :	result = 16'd6;
         64600    :	result = 16'd6;
         64601    :	result = 16'd6;
         64602    :	result = 16'd6;
         64603    :	result = 16'd6;
         64604    :	result = 16'd6;
         64605    :	result = 16'd6;
         64606    :	result = 16'd6;
         64607    :	result = 16'd6;
         64608    :	result = 16'd6;
         64609    :	result = 16'd6;
         64610    :	result = 16'd6;
         64611    :	result = 16'd6;
         64612    :	result = 16'd6;
         64613    :	result = 16'd6;
         64614    :	result = 16'd6;
         64615    :	result = 16'd6;
         64616    :	result = 16'd6;
         64617    :	result = 16'd6;
         64618    :	result = 16'd6;
         64619    :	result = 16'd6;
         64620    :	result = 16'd6;
         64621    :	result = 16'd7;
         64622    :	result = 16'd7;
         64623    :	result = 16'd7;
         64624    :	result = 16'd7;
         64625    :	result = 16'd7;
         64626    :	result = 16'd7;
         64627    :	result = 16'd7;
         64628    :	result = 16'd7;
         64629    :	result = 16'd7;
         64630    :	result = 16'd7;
         64631    :	result = 16'd7;
         64632    :	result = 16'd7;
         64633    :	result = 16'd7;
         64634    :	result = 16'd7;
         64635    :	result = 16'd7;
         64636    :	result = 16'd7;
         64637    :	result = 16'd7;
         64638    :	result = 16'd7;
         64639    :	result = 16'd7;
         64640    :	result = 16'd7;
         64641    :	result = 16'd7;
         64642    :	result = 16'd7;
         64643    :	result = 16'd7;
         64644    :	result = 16'd7;
         64645    :	result = 16'd7;
         64646    :	result = 16'd7;
         64647    :	result = 16'd7;
         64648    :	result = 16'd7;
         64649    :	result = 16'd7;
         64650    :	result = 16'd7;
         64651    :	result = 16'd7;
         64652    :	result = 16'd7;
         64653    :	result = 16'd7;
         64654    :	result = 16'd7;
         64655    :	result = 16'd7;
         64656    :	result = 16'd8;
         64657    :	result = 16'd8;
         64658    :	result = 16'd8;
         64659    :	result = 16'd8;
         64660    :	result = 16'd8;
         64661    :	result = 16'd8;
         64662    :	result = 16'd8;
         64663    :	result = 16'd8;
         64664    :	result = 16'd8;
         64665    :	result = 16'd8;
         64666    :	result = 16'd8;
         64667    :	result = 16'd8;
         64668    :	result = 16'd8;
         64669    :	result = 16'd8;
         64670    :	result = 16'd8;
         64671    :	result = 16'd8;
         64672    :	result = 16'd8;
         64673    :	result = 16'd8;
         64674    :	result = 16'd8;
         64675    :	result = 16'd8;
         64676    :	result = 16'd8;
         64677    :	result = 16'd8;
         64678    :	result = 16'd8;
         64679    :	result = 16'd8;
         64680    :	result = 16'd8;
         64681    :	result = 16'd8;
         64682    :	result = 16'd8;
         64683    :	result = 16'd8;
         64684    :	result = 16'd8;
         64685    :	result = 16'd8;
         64686    :	result = 16'd8;
         64687    :	result = 16'd8;
         64688    :	result = 16'd9;
         64689    :	result = 16'd9;
         64690    :	result = 16'd9;
         64691    :	result = 16'd9;
         64692    :	result = 16'd9;
         64693    :	result = 16'd9;
         64694    :	result = 16'd9;
         64695    :	result = 16'd9;
         64696    :	result = 16'd9;
         64697    :	result = 16'd9;
         64698    :	result = 16'd9;
         64699    :	result = 16'd9;
         64700    :	result = 16'd9;
         64701    :	result = 16'd9;
         64702    :	result = 16'd9;
         64703    :	result = 16'd9;
         64704    :	result = 16'd9;
         64705    :	result = 16'd9;
         64706    :	result = 16'd9;
         64707    :	result = 16'd9;
         64708    :	result = 16'd9;
         64709    :	result = 16'd9;
         64710    :	result = 16'd9;
         64711    :	result = 16'd9;
         64712    :	result = 16'd9;
         64713    :	result = 16'd9;
         64714    :	result = 16'd9;
         64715    :	result = 16'd9;
         64716    :	result = 16'd10;
         64717    :	result = 16'd10;
         64718    :	result = 16'd10;
         64719    :	result = 16'd10;
         64720    :	result = 16'd10;
         64721    :	result = 16'd10;
         64722    :	result = 16'd10;
         64723    :	result = 16'd10;
         64724    :	result = 16'd10;
         64725    :	result = 16'd10;
         64726    :	result = 16'd10;
         64727    :	result = 16'd10;
         64728    :	result = 16'd10;
         64729    :	result = 16'd10;
         64730    :	result = 16'd10;
         64731    :	result = 16'd10;
         64732    :	result = 16'd10;
         64733    :	result = 16'd10;
         64734    :	result = 16'd10;
         64735    :	result = 16'd10;
         64736    :	result = 16'd10;
         64737    :	result = 16'd10;
         64738    :	result = 16'd10;
         64739    :	result = 16'd10;
         64740    :	result = 16'd10;
         64741    :	result = 16'd11;
         64742    :	result = 16'd11;
         64743    :	result = 16'd11;
         64744    :	result = 16'd11;
         64745    :	result = 16'd11;
         64746    :	result = 16'd11;
         64747    :	result = 16'd11;
         64748    :	result = 16'd11;
         64749    :	result = 16'd11;
         64750    :	result = 16'd11;
         64751    :	result = 16'd11;
         64752    :	result = 16'd11;
         64753    :	result = 16'd11;
         64754    :	result = 16'd11;
         64755    :	result = 16'd11;
         64756    :	result = 16'd11;
         64757    :	result = 16'd11;
         64758    :	result = 16'd11;
         64759    :	result = 16'd11;
         64760    :	result = 16'd11;
         64761    :	result = 16'd11;
         64762    :	result = 16'd11;
         64763    :	result = 16'd11;
         64764    :	result = 16'd12;
         64765    :	result = 16'd12;
         64766    :	result = 16'd12;
         64767    :	result = 16'd12;
         64768    :	result = 16'd12;
         64769    :	result = 16'd12;
         64770    :	result = 16'd12;
         64771    :	result = 16'd12;
         64772    :	result = 16'd12;
         64773    :	result = 16'd12;
         64774    :	result = 16'd12;
         64775    :	result = 16'd12;
         64776    :	result = 16'd12;
         64777    :	result = 16'd12;
         64778    :	result = 16'd12;
         64779    :	result = 16'd12;
         64780    :	result = 16'd12;
         64781    :	result = 16'd12;
         64782    :	result = 16'd12;
         64783    :	result = 16'd12;
         64784    :	result = 16'd12;
         64785    :	result = 16'd12;
         64786    :	result = 16'd13;
         64787    :	result = 16'd13;
         64788    :	result = 16'd13;
         64789    :	result = 16'd13;
         64790    :	result = 16'd13;
         64791    :	result = 16'd13;
         64792    :	result = 16'd13;
         64793    :	result = 16'd13;
         64794    :	result = 16'd13;
         64795    :	result = 16'd13;
         64796    :	result = 16'd13;
         64797    :	result = 16'd13;
         64798    :	result = 16'd13;
         64799    :	result = 16'd13;
         64800    :	result = 16'd13;
         64801    :	result = 16'd13;
         64802    :	result = 16'd13;
         64803    :	result = 16'd13;
         64804    :	result = 16'd13;
         64805    :	result = 16'd13;
         64806    :	result = 16'd14;
         64807    :	result = 16'd14;
         64808    :	result = 16'd14;
         64809    :	result = 16'd14;
         64810    :	result = 16'd14;
         64811    :	result = 16'd14;
         64812    :	result = 16'd14;
         64813    :	result = 16'd14;
         64814    :	result = 16'd14;
         64815    :	result = 16'd14;
         64816    :	result = 16'd14;
         64817    :	result = 16'd14;
         64818    :	result = 16'd14;
         64819    :	result = 16'd14;
         64820    :	result = 16'd14;
         64821    :	result = 16'd14;
         64822    :	result = 16'd14;
         64823    :	result = 16'd14;
         64824    :	result = 16'd14;
         64825    :	result = 16'd15;
         64826    :	result = 16'd15;
         64827    :	result = 16'd15;
         64828    :	result = 16'd15;
         64829    :	result = 16'd15;
         64830    :	result = 16'd15;
         64831    :	result = 16'd15;
         64832    :	result = 16'd15;
         64833    :	result = 16'd15;
         64834    :	result = 16'd15;
         64835    :	result = 16'd15;
         64836    :	result = 16'd15;
         64837    :	result = 16'd15;
         64838    :	result = 16'd15;
         64839    :	result = 16'd15;
         64840    :	result = 16'd15;
         64841    :	result = 16'd15;
         64842    :	result = 16'd16;
         64843    :	result = 16'd16;
         64844    :	result = 16'd16;
         64845    :	result = 16'd16;
         64846    :	result = 16'd16;
         64847    :	result = 16'd16;
         64848    :	result = 16'd16;
         64849    :	result = 16'd16;
         64850    :	result = 16'd16;
         64851    :	result = 16'd16;
         64852    :	result = 16'd16;
         64853    :	result = 16'd16;
         64854    :	result = 16'd16;
         64855    :	result = 16'd16;
         64856    :	result = 16'd16;
         64857    :	result = 16'd16;
         64858    :	result = 16'd16;
         64859    :	result = 16'd17;
         64860    :	result = 16'd17;
         64861    :	result = 16'd17;
         64862    :	result = 16'd17;
         64863    :	result = 16'd17;
         64864    :	result = 16'd17;
         64865    :	result = 16'd17;
         64866    :	result = 16'd17;
         64867    :	result = 16'd17;
         64868    :	result = 16'd17;
         64869    :	result = 16'd17;
         64870    :	result = 16'd17;
         64871    :	result = 16'd17;
         64872    :	result = 16'd17;
         64873    :	result = 16'd17;
         64874    :	result = 16'd17;
         64875    :	result = 16'd18;
         64876    :	result = 16'd18;
         64877    :	result = 16'd18;
         64878    :	result = 16'd18;
         64879    :	result = 16'd18;
         64880    :	result = 16'd18;
         64881    :	result = 16'd18;
         64882    :	result = 16'd18;
         64883    :	result = 16'd18;
         64884    :	result = 16'd18;
         64885    :	result = 16'd18;
         64886    :	result = 16'd18;
         64887    :	result = 16'd18;
         64888    :	result = 16'd18;
         64889    :	result = 16'd19;
         64890    :	result = 16'd19;
         64891    :	result = 16'd19;
         64892    :	result = 16'd19;
         64893    :	result = 16'd19;
         64894    :	result = 16'd19;
         64895    :	result = 16'd19;
         64896    :	result = 16'd19;
         64897    :	result = 16'd19;
         64898    :	result = 16'd19;
         64899    :	result = 16'd19;
         64900    :	result = 16'd19;
         64901    :	result = 16'd19;
         64902    :	result = 16'd19;
         64903    :	result = 16'd19;
         64904    :	result = 16'd20;
         64905    :	result = 16'd20;
         64906    :	result = 16'd20;
         64907    :	result = 16'd20;
         64908    :	result = 16'd20;
         64909    :	result = 16'd20;
         64910    :	result = 16'd20;
         64911    :	result = 16'd20;
         64912    :	result = 16'd20;
         64913    :	result = 16'd20;
         64914    :	result = 16'd20;
         64915    :	result = 16'd20;
         64916    :	result = 16'd20;
         64917    :	result = 16'd21;
         64918    :	result = 16'd21;
         64919    :	result = 16'd21;
         64920    :	result = 16'd21;
         64921    :	result = 16'd21;
         64922    :	result = 16'd21;
         64923    :	result = 16'd21;
         64924    :	result = 16'd21;
         64925    :	result = 16'd21;
         64926    :	result = 16'd21;
         64927    :	result = 16'd21;
         64928    :	result = 16'd21;
         64929    :	result = 16'd21;
         64930    :	result = 16'd22;
         64931    :	result = 16'd22;
         64932    :	result = 16'd22;
         64933    :	result = 16'd22;
         64934    :	result = 16'd22;
         64935    :	result = 16'd22;
         64936    :	result = 16'd22;
         64937    :	result = 16'd22;
         64938    :	result = 16'd22;
         64939    :	result = 16'd22;
         64940    :	result = 16'd22;
         64941    :	result = 16'd22;
         64942    :	result = 16'd22;
         64943    :	result = 16'd23;
         64944    :	result = 16'd23;
         64945    :	result = 16'd23;
         64946    :	result = 16'd23;
         64947    :	result = 16'd23;
         64948    :	result = 16'd23;
         64949    :	result = 16'd23;
         64950    :	result = 16'd23;
         64951    :	result = 16'd23;
         64952    :	result = 16'd23;
         64953    :	result = 16'd23;
         64954    :	result = 16'd23;
         64955    :	result = 16'd24;
         64956    :	result = 16'd24;
         64957    :	result = 16'd24;
         64958    :	result = 16'd24;
         64959    :	result = 16'd24;
         64960    :	result = 16'd24;
         64961    :	result = 16'd24;
         64962    :	result = 16'd24;
         64963    :	result = 16'd24;
         64964    :	result = 16'd24;
         64965    :	result = 16'd24;
         64966    :	result = 16'd25;
         64967    :	result = 16'd25;
         64968    :	result = 16'd25;
         64969    :	result = 16'd25;
         64970    :	result = 16'd25;
         64971    :	result = 16'd25;
         64972    :	result = 16'd25;
         64973    :	result = 16'd25;
         64974    :	result = 16'd25;
         64975    :	result = 16'd25;
         64976    :	result = 16'd25;
         64977    :	result = 16'd26;
         64978    :	result = 16'd26;
         64979    :	result = 16'd26;
         64980    :	result = 16'd26;
         64981    :	result = 16'd26;
         64982    :	result = 16'd26;
         64983    :	result = 16'd26;
         64984    :	result = 16'd26;
         64985    :	result = 16'd26;
         64986    :	result = 16'd26;
         64987    :	result = 16'd26;
         64988    :	result = 16'd27;
         64989    :	result = 16'd27;
         64990    :	result = 16'd27;
         64991    :	result = 16'd27;
         64992    :	result = 16'd27;
         64993    :	result = 16'd27;
         64994    :	result = 16'd27;
         64995    :	result = 16'd27;
         64996    :	result = 16'd27;
         64997    :	result = 16'd27;
         64998    :	result = 16'd27;
         64999    :	result = 16'd28;
         65000    :	result = 16'd28;
         65001    :	result = 16'd28;
         65002    :	result = 16'd28;
         65003    :	result = 16'd28;
         65004    :	result = 16'd28;
         65005    :	result = 16'd28;
         65006    :	result = 16'd28;
         65007    :	result = 16'd28;
         65008    :	result = 16'd28;
         65009    :	result = 16'd29;
         65010    :	result = 16'd29;
         65011    :	result = 16'd29;
         65012    :	result = 16'd29;
         65013    :	result = 16'd29;
         65014    :	result = 16'd29;
         65015    :	result = 16'd29;
         65016    :	result = 16'd29;
         65017    :	result = 16'd29;
         65018    :	result = 16'd29;
         65019    :	result = 16'd30;
         65020    :	result = 16'd30;
         65021    :	result = 16'd30;
         65022    :	result = 16'd30;
         65023    :	result = 16'd30;
         65024    :	result = 16'd30;
         65025    :	result = 16'd30;
         65026    :	result = 16'd30;
         65027    :	result = 16'd30;
         65028    :	result = 16'd31;
         65029    :	result = 16'd31;
         65030    :	result = 16'd31;
         65031    :	result = 16'd31;
         65032    :	result = 16'd31;
         65033    :	result = 16'd31;
         65034    :	result = 16'd31;
         65035    :	result = 16'd31;
         65036    :	result = 16'd31;
         65037    :	result = 16'd32;
         65038    :	result = 16'd32;
         65039    :	result = 16'd32;
         65040    :	result = 16'd32;
         65041    :	result = 16'd32;
         65042    :	result = 16'd32;
         65043    :	result = 16'd32;
         65044    :	result = 16'd32;
         65045    :	result = 16'd32;
         65046    :	result = 16'd33;
         65047    :	result = 16'd33;
         65048    :	result = 16'd33;
         65049    :	result = 16'd33;
         65050    :	result = 16'd33;
         65051    :	result = 16'd33;
         65052    :	result = 16'd33;
         65053    :	result = 16'd33;
         65054    :	result = 16'd33;
         65055    :	result = 16'd34;
         65056    :	result = 16'd34;
         65057    :	result = 16'd34;
         65058    :	result = 16'd34;
         65059    :	result = 16'd34;
         65060    :	result = 16'd34;
         65061    :	result = 16'd34;
         65062    :	result = 16'd34;
         65063    :	result = 16'd34;
         65064    :	result = 16'd35;
         65065    :	result = 16'd35;
         65066    :	result = 16'd35;
         65067    :	result = 16'd35;
         65068    :	result = 16'd35;
         65069    :	result = 16'd35;
         65070    :	result = 16'd35;
         65071    :	result = 16'd35;
         65072    :	result = 16'd36;
         65073    :	result = 16'd36;
         65074    :	result = 16'd36;
         65075    :	result = 16'd36;
         65076    :	result = 16'd36;
         65077    :	result = 16'd36;
         65078    :	result = 16'd36;
         65079    :	result = 16'd36;
         65080    :	result = 16'd37;
         65081    :	result = 16'd37;
         65082    :	result = 16'd37;
         65083    :	result = 16'd37;
         65084    :	result = 16'd37;
         65085    :	result = 16'd37;
         65086    :	result = 16'd37;
         65087    :	result = 16'd37;
         65088    :	result = 16'd38;
         65089    :	result = 16'd38;
         65090    :	result = 16'd38;
         65091    :	result = 16'd38;
         65092    :	result = 16'd38;
         65093    :	result = 16'd38;
         65094    :	result = 16'd38;
         65095    :	result = 16'd38;
         65096    :	result = 16'd39;
         65097    :	result = 16'd39;
         65098    :	result = 16'd39;
         65099    :	result = 16'd39;
         65100    :	result = 16'd39;
         65101    :	result = 16'd39;
         65102    :	result = 16'd39;
         65103    :	result = 16'd39;
         65104    :	result = 16'd40;
         65105    :	result = 16'd40;
         65106    :	result = 16'd40;
         65107    :	result = 16'd40;
         65108    :	result = 16'd40;
         65109    :	result = 16'd40;
         65110    :	result = 16'd40;
         65111    :	result = 16'd41;
         65112    :	result = 16'd41;
         65113    :	result = 16'd41;
         65114    :	result = 16'd41;
         65115    :	result = 16'd41;
         65116    :	result = 16'd41;
         65117    :	result = 16'd41;
         65118    :	result = 16'd41;
         65119    :	result = 16'd42;
         65120    :	result = 16'd42;
         65121    :	result = 16'd42;
         65122    :	result = 16'd42;
         65123    :	result = 16'd42;
         65124    :	result = 16'd42;
         65125    :	result = 16'd42;
         65126    :	result = 16'd43;
         65127    :	result = 16'd43;
         65128    :	result = 16'd43;
         65129    :	result = 16'd43;
         65130    :	result = 16'd43;
         65131    :	result = 16'd43;
         65132    :	result = 16'd43;
         65133    :	result = 16'd44;
         65134    :	result = 16'd44;
         65135    :	result = 16'd44;
         65136    :	result = 16'd44;
         65137    :	result = 16'd44;
         65138    :	result = 16'd44;
         65139    :	result = 16'd44;
         65140    :	result = 16'd45;
         65141    :	result = 16'd45;
         65142    :	result = 16'd45;
         65143    :	result = 16'd45;
         65144    :	result = 16'd45;
         65145    :	result = 16'd45;
         65146    :	result = 16'd45;
         65147    :	result = 16'd46;
         65148    :	result = 16'd46;
         65149    :	result = 16'd46;
         65150    :	result = 16'd46;
         65151    :	result = 16'd46;
         65152    :	result = 16'd46;
         65153    :	result = 16'd46;
         65154    :	result = 16'd47;
         65155    :	result = 16'd47;
         65156    :	result = 16'd47;
         65157    :	result = 16'd47;
         65158    :	result = 16'd47;
         65159    :	result = 16'd47;
         65160    :	result = 16'd48;
         65161    :	result = 16'd48;
         65162    :	result = 16'd48;
         65163    :	result = 16'd48;
         65164    :	result = 16'd48;
         65165    :	result = 16'd48;
         65166    :	result = 16'd48;
         65167    :	result = 16'd49;
         65168    :	result = 16'd49;
         65169    :	result = 16'd49;
         65170    :	result = 16'd49;
         65171    :	result = 16'd49;
         65172    :	result = 16'd49;
         65173    :	result = 16'd50;
         65174    :	result = 16'd50;
         65175    :	result = 16'd50;
         65176    :	result = 16'd50;
         65177    :	result = 16'd50;
         65178    :	result = 16'd50;
         65179    :	result = 16'd51;
         65180    :	result = 16'd51;
         65181    :	result = 16'd51;
         65182    :	result = 16'd51;
         65183    :	result = 16'd51;
         65184    :	result = 16'd51;
         65185    :	result = 16'd51;
         65186    :	result = 16'd52;
         65187    :	result = 16'd52;
         65188    :	result = 16'd52;
         65189    :	result = 16'd52;
         65190    :	result = 16'd52;
         65191    :	result = 16'd52;
         65192    :	result = 16'd53;
         65193    :	result = 16'd53;
         65194    :	result = 16'd53;
         65195    :	result = 16'd53;
         65196    :	result = 16'd53;
         65197    :	result = 16'd53;
         65198    :	result = 16'd54;
         65199    :	result = 16'd54;
         65200    :	result = 16'd54;
         65201    :	result = 16'd54;
         65202    :	result = 16'd54;
         65203    :	result = 16'd54;
         65204    :	result = 16'd55;
         65205    :	result = 16'd55;
         65206    :	result = 16'd55;
         65207    :	result = 16'd55;
         65208    :	result = 16'd55;
         65209    :	result = 16'd55;
         65210    :	result = 16'd56;
         65211    :	result = 16'd56;
         65212    :	result = 16'd56;
         65213    :	result = 16'd56;
         65214    :	result = 16'd56;
         65215    :	result = 16'd57;
         65216    :	result = 16'd57;
         65217    :	result = 16'd57;
         65218    :	result = 16'd57;
         65219    :	result = 16'd57;
         65220    :	result = 16'd57;
         65221    :	result = 16'd58;
         65222    :	result = 16'd58;
         65223    :	result = 16'd58;
         65224    :	result = 16'd58;
         65225    :	result = 16'd58;
         65226    :	result = 16'd58;
         65227    :	result = 16'd59;
         65228    :	result = 16'd59;
         65229    :	result = 16'd59;
         65230    :	result = 16'd59;
         65231    :	result = 16'd59;
         65232    :	result = 16'd60;
         65233    :	result = 16'd60;
         65234    :	result = 16'd60;
         65235    :	result = 16'd60;
         65236    :	result = 16'd60;
         65237    :	result = 16'd60;
         65238    :	result = 16'd61;
         65239    :	result = 16'd61;
         65240    :	result = 16'd61;
         65241    :	result = 16'd61;
         65242    :	result = 16'd61;
         65243    :	result = 16'd62;
         65244    :	result = 16'd62;
         65245    :	result = 16'd62;
         65246    :	result = 16'd62;
         65247    :	result = 16'd62;
         65248    :	result = 16'd62;
         65249    :	result = 16'd63;
         65250    :	result = 16'd63;
         65251    :	result = 16'd63;
         65252    :	result = 16'd63;
         65253    :	result = 16'd63;
         65254    :	result = 16'd64;
         65255    :	result = 16'd64;
         65256    :	result = 16'd64;
         65257    :	result = 16'd64;
         65258    :	result = 16'd64;
         65259    :	result = 16'd64;
         65260    :	result = 16'd65;
         65261    :	result = 16'd65;
         65262    :	result = 16'd65;
         65263    :	result = 16'd65;
         65264    :	result = 16'd65;
         65265    :	result = 16'd66;
         65266    :	result = 16'd66;
         65267    :	result = 16'd66;
         65268    :	result = 16'd66;
         65269    :	result = 16'd66;
         65270    :	result = 16'd67;
         65271    :	result = 16'd67;
         65272    :	result = 16'd67;
         65273    :	result = 16'd67;
         65274    :	result = 16'd67;
         65275    :	result = 16'd68;
         65276    :	result = 16'd68;
         65277    :	result = 16'd68;
         65278    :	result = 16'd68;
         65279    :	result = 16'd68;
         65280    :	result = 16'd69;
         65281    :	result = 16'd69;
         65282    :	result = 16'd69;
         65283    :	result = 16'd69;
         65284    :	result = 16'd69;
         65285    :	result = 16'd70;
         65286    :	result = 16'd70;
         65287    :	result = 16'd70;
         65288    :	result = 16'd70;
         65289    :	result = 16'd70;
         65290    :	result = 16'd71;
         65291    :	result = 16'd71;
         65292    :	result = 16'd71;
         65293    :	result = 16'd71;
         65294    :	result = 16'd71;
         65295    :	result = 16'd72;
         65296    :	result = 16'd72;
         65297    :	result = 16'd72;
         65298    :	result = 16'd72;
         65299    :	result = 16'd72;
         65300    :	result = 16'd73;
         65301    :	result = 16'd73;
         65302    :	result = 16'd73;
         65303    :	result = 16'd73;
         65304    :	result = 16'd73;
         65305    :	result = 16'd74;
         65306    :	result = 16'd74;
         65307    :	result = 16'd74;
         65308    :	result = 16'd74;
         65309    :	result = 16'd74;
         65310    :	result = 16'd75;
         65311    :	result = 16'd75;
         65312    :	result = 16'd75;
         65313    :	result = 16'd75;
         65314    :	result = 16'd75;
         65315    :	result = 16'd76;
         65316    :	result = 16'd76;
         65317    :	result = 16'd76;
         65318    :	result = 16'd76;
         65319    :	result = 16'd76;
         65320    :	result = 16'd77;
         65321    :	result = 16'd77;
         65322    :	result = 16'd77;
         65323    :	result = 16'd77;
         65324    :	result = 16'd78;
         65325    :	result = 16'd78;
         65326    :	result = 16'd78;
         65327    :	result = 16'd78;
         65328    :	result = 16'd78;
         65329    :	result = 16'd79;
         65330    :	result = 16'd79;
         65331    :	result = 16'd79;
         65332    :	result = 16'd79;
         65333    :	result = 16'd79;
         65334    :	result = 16'd80;
         65335    :	result = 16'd80;
         65336    :	result = 16'd80;
         65337    :	result = 16'd80;
         65338    :	result = 16'd81;
         65339    :	result = 16'd81;
         65340    :	result = 16'd81;
         65341    :	result = 16'd81;
         65342    :	result = 16'd81;
         65343    :	result = 16'd82;
         65344    :	result = 16'd82;
         65345    :	result = 16'd82;
         65346    :	result = 16'd82;
         65347    :	result = 16'd83;
         65348    :	result = 16'd83;
         65349    :	result = 16'd83;
         65350    :	result = 16'd83;
         65351    :	result = 16'd83;
         65352    :	result = 16'd84;
         65353    :	result = 16'd84;
         65354    :	result = 16'd84;
         65355    :	result = 16'd84;
         65356    :	result = 16'd84;
         65357    :	result = 16'd85;
         65358    :	result = 16'd85;
         65359    :	result = 16'd85;
         65360    :	result = 16'd85;
         65361    :	result = 16'd86;
         65362    :	result = 16'd86;
         65363    :	result = 16'd86;
         65364    :	result = 16'd86;
         65365    :	result = 16'd86;
         65366    :	result = 16'd87;
         65367    :	result = 16'd87;
         65368    :	result = 16'd87;
         65369    :	result = 16'd87;
         65370    :	result = 16'd88;
         65371    :	result = 16'd88;
         65372    :	result = 16'd88;
         65373    :	result = 16'd88;
         65374    :	result = 16'd89;
         65375    :	result = 16'd89;
         65376    :	result = 16'd89;
         65377    :	result = 16'd89;
         65378    :	result = 16'd89;
         65379    :	result = 16'd90;
         65380    :	result = 16'd90;
         65381    :	result = 16'd90;
         65382    :	result = 16'd90;
         65383    :	result = 16'd91;
         65384    :	result = 16'd91;
         65385    :	result = 16'd91;
         65386    :	result = 16'd91;
         65387    :	result = 16'd91;
         65388    :	result = 16'd92;
         65389    :	result = 16'd92;
         65390    :	result = 16'd92;
         65391    :	result = 16'd92;
         65392    :	result = 16'd93;
         65393    :	result = 16'd93;
         65394    :	result = 16'd93;
         65395    :	result = 16'd93;
         65396    :	result = 16'd94;
         65397    :	result = 16'd94;
         65398    :	result = 16'd94;
         65399    :	result = 16'd94;
         65400    :	result = 16'd95;
         65401    :	result = 16'd95;
         65402    :	result = 16'd95;
         65403    :	result = 16'd95;
         65404    :	result = 16'd95;
         65405    :	result = 16'd96;
         65406    :	result = 16'd96;
         65407    :	result = 16'd96;
         65408    :	result = 16'd96;
         65409    :	result = 16'd97;
         65410    :	result = 16'd97;
         65411    :	result = 16'd97;
         65412    :	result = 16'd97;
         65413    :	result = 16'd98;
         65414    :	result = 16'd98;
         65415    :	result = 16'd98;
         65416    :	result = 16'd98;
         65417    :	result = 16'd99;
         65418    :	result = 16'd99;
         65419    :	result = 16'd99;
         65420    :	result = 16'd99;
         65421    :	result = 16'd99;
         65422    :	result = 16'd100;
         65423    :	result = 16'd100;
         65424    :	result = 16'd100;
         65425    :	result = 16'd100;
         65426    :	result = 16'd101;
         65427    :	result = 16'd101;
         65428    :	result = 16'd101;
         65429    :	result = 16'd101;
         65430    :	result = 16'd102;
         65431    :	result = 16'd102;
         65432    :	result = 16'd102;
         65433    :	result = 16'd102;
         65434    :	result = 16'd103;
         65435    :	result = 16'd103;
         65436    :	result = 16'd103;
         65437    :	result = 16'd103;
         65438    :	result = 16'd104;
         65439    :	result = 16'd104;
         65440    :	result = 16'd104;
         65441    :	result = 16'd104;
         65442    :	result = 16'd105;
         65443    :	result = 16'd105;
         65444    :	result = 16'd105;
         65445    :	result = 16'd105;
         65446    :	result = 16'd105;
         65447    :	result = 16'd106;
         65448    :	result = 16'd106;
         65449    :	result = 16'd106;
         65450    :	result = 16'd106;
         65451    :	result = 16'd107;
         65452    :	result = 16'd107;
         65453    :	result = 16'd107;
         65454    :	result = 16'd107;
         65455    :	result = 16'd108;
         65456    :	result = 16'd108;
         65457    :	result = 16'd108;
         65458    :	result = 16'd108;
         65459    :	result = 16'd109;
         65460    :	result = 16'd109;
         65461    :	result = 16'd109;
         65462    :	result = 16'd109;
         65463    :	result = 16'd110;
         65464    :	result = 16'd110;
         65465    :	result = 16'd110;
         65466    :	result = 16'd110;
         65467    :	result = 16'd111;
         65468    :	result = 16'd111;
         65469    :	result = 16'd111;
         65470    :	result = 16'd111;
         65471    :	result = 16'd112;
         65472    :	result = 16'd112;
         65473    :	result = 16'd112;
         65474    :	result = 16'd112;
         65475    :	result = 16'd113;
         65476    :	result = 16'd113;
         65477    :	result = 16'd113;
         65478    :	result = 16'd113;
         65479    :	result = 16'd114;
         65480    :	result = 16'd114;
         65481    :	result = 16'd114;
         65482    :	result = 16'd114;
         65483    :	result = 16'd115;
         65484    :	result = 16'd115;
         65485    :	result = 16'd115;
         65486    :	result = 16'd115;
         65487    :	result = 16'd116;
         65488    :	result = 16'd116;
         65489    :	result = 16'd116;
         65490    :	result = 16'd116;
         65491    :	result = 16'd117;
         65492    :	result = 16'd117;
         65493    :	result = 16'd117;
         65494    :	result = 16'd117;
         65495    :	result = 16'd118;
         65496    :	result = 16'd118;
         65497    :	result = 16'd118;
         65498    :	result = 16'd118;
         65499    :	result = 16'd119;
         65500    :	result = 16'd119;
         65501    :	result = 16'd119;
         65502    :	result = 16'd119;
         65503    :	result = 16'd120;
         65504    :	result = 16'd120;
         65505    :	result = 16'd120;
         65506    :	result = 16'd120;
         65507    :	result = 16'd121;
         65508    :	result = 16'd121;
         65509    :	result = 16'd121;
         65510    :	result = 16'd121;
         65511    :	result = 16'd122;
         65512    :	result = 16'd122;
         65513    :	result = 16'd122;
         65514    :	result = 16'd122;
         65515    :	result = 16'd123;
         65516    :	result = 16'd123;
         65517    :	result = 16'd123;
         65518    :	result = 16'd123;
         65519    :	result = 16'd124;
         65520    :	result = 16'd124;
         65521    :	result = 16'd124;
         65522    :	result = 16'd124;
         65523    :	result = 16'd125;
         65524    :	result = 16'd125;
         65525    :	result = 16'd125;
         65526    :	result = 16'd125;
         65527    :	result = 16'd126;
         65528    :	result = 16'd126;
         65529    :	result = 16'd126;
         65530    :	result = 16'd126;
         65531    :	result = 16'd127;
         65532    :	result = 16'd127;
         65533    :	result = 16'd127;
         65534    :	result = 16'd127;
         65535    :	result = 16'd128;
         0        :	result = 16'd128;
         1        :	result = 16'd128;
         2        :	result = 16'd128;
         3        :	result = 16'd128;
         4        :	result = 16'd129;
         5        :	result = 16'd129;
         6        :	result = 16'd129;
         7        :	result = 16'd129;
         8        :	result = 16'd130;
         9        :	result = 16'd130;
         10       :	result = 16'd130;
         11       :	result = 16'd130;
         12       :	result = 16'd131;
         13       :	result = 16'd131;
         14       :	result = 16'd131;
         15       :	result = 16'd131;
         16       :	result = 16'd132;
         17       :	result = 16'd132;
         18       :	result = 16'd132;
         19       :	result = 16'd132;
         20       :	result = 16'd133;
         21       :	result = 16'd133;
         22       :	result = 16'd133;
         23       :	result = 16'd133;
         24       :	result = 16'd134;
         25       :	result = 16'd134;
         26       :	result = 16'd134;
         27       :	result = 16'd134;
         28       :	result = 16'd135;
         29       :	result = 16'd135;
         30       :	result = 16'd135;
         31       :	result = 16'd135;
         32       :	result = 16'd136;
         33       :	result = 16'd136;
         34       :	result = 16'd136;
         35       :	result = 16'd136;
         36       :	result = 16'd137;
         37       :	result = 16'd137;
         38       :	result = 16'd137;
         39       :	result = 16'd137;
         40       :	result = 16'd138;
         41       :	result = 16'd138;
         42       :	result = 16'd138;
         43       :	result = 16'd138;
         44       :	result = 16'd139;
         45       :	result = 16'd139;
         46       :	result = 16'd139;
         47       :	result = 16'd139;
         48       :	result = 16'd140;
         49       :	result = 16'd140;
         50       :	result = 16'd140;
         51       :	result = 16'd140;
         52       :	result = 16'd141;
         53       :	result = 16'd141;
         54       :	result = 16'd141;
         55       :	result = 16'd141;
         56       :	result = 16'd142;
         57       :	result = 16'd142;
         58       :	result = 16'd142;
         59       :	result = 16'd142;
         60       :	result = 16'd143;
         61       :	result = 16'd143;
         62       :	result = 16'd143;
         63       :	result = 16'd143;
         64       :	result = 16'd144;
         65       :	result = 16'd144;
         66       :	result = 16'd144;
         67       :	result = 16'd144;
         68       :	result = 16'd145;
         69       :	result = 16'd145;
         70       :	result = 16'd145;
         71       :	result = 16'd145;
         72       :	result = 16'd146;
         73       :	result = 16'd146;
         74       :	result = 16'd146;
         75       :	result = 16'd146;
         76       :	result = 16'd147;
         77       :	result = 16'd147;
         78       :	result = 16'd147;
         79       :	result = 16'd147;
         80       :	result = 16'd148;
         81       :	result = 16'd148;
         82       :	result = 16'd148;
         83       :	result = 16'd148;
         84       :	result = 16'd149;
         85       :	result = 16'd149;
         86       :	result = 16'd149;
         87       :	result = 16'd149;
         88       :	result = 16'd150;
         89       :	result = 16'd150;
         90       :	result = 16'd150;
         91       :	result = 16'd150;
         92       :	result = 16'd150;
         93       :	result = 16'd151;
         94       :	result = 16'd151;
         95       :	result = 16'd151;
         96       :	result = 16'd151;
         97       :	result = 16'd152;
         98       :	result = 16'd152;
         99       :	result = 16'd152;
         100      :	result = 16'd152;
         101      :	result = 16'd153;
         102      :	result = 16'd153;
         103      :	result = 16'd153;
         104      :	result = 16'd153;
         105      :	result = 16'd154;
         106      :	result = 16'd154;
         107      :	result = 16'd154;
         108      :	result = 16'd154;
         109      :	result = 16'd155;
         110      :	result = 16'd155;
         111      :	result = 16'd155;
         112      :	result = 16'd155;
         113      :	result = 16'd156;
         114      :	result = 16'd156;
         115      :	result = 16'd156;
         116      :	result = 16'd156;
         117      :	result = 16'd156;
         118      :	result = 16'd157;
         119      :	result = 16'd157;
         120      :	result = 16'd157;
         121      :	result = 16'd157;
         122      :	result = 16'd158;
         123      :	result = 16'd158;
         124      :	result = 16'd158;
         125      :	result = 16'd158;
         126      :	result = 16'd159;
         127      :	result = 16'd159;
         128      :	result = 16'd159;
         129      :	result = 16'd159;
         130      :	result = 16'd160;
         131      :	result = 16'd160;
         132      :	result = 16'd160;
         133      :	result = 16'd160;
         134      :	result = 16'd160;
         135      :	result = 16'd161;
         136      :	result = 16'd161;
         137      :	result = 16'd161;
         138      :	result = 16'd161;
         139      :	result = 16'd162;
         140      :	result = 16'd162;
         141      :	result = 16'd162;
         142      :	result = 16'd162;
         143      :	result = 16'd163;
         144      :	result = 16'd163;
         145      :	result = 16'd163;
         146      :	result = 16'd163;
         147      :	result = 16'd164;
         148      :	result = 16'd164;
         149      :	result = 16'd164;
         150      :	result = 16'd164;
         151      :	result = 16'd164;
         152      :	result = 16'd165;
         153      :	result = 16'd165;
         154      :	result = 16'd165;
         155      :	result = 16'd165;
         156      :	result = 16'd166;
         157      :	result = 16'd166;
         158      :	result = 16'd166;
         159      :	result = 16'd166;
         160      :	result = 16'd166;
         161      :	result = 16'd167;
         162      :	result = 16'd167;
         163      :	result = 16'd167;
         164      :	result = 16'd167;
         165      :	result = 16'd168;
         166      :	result = 16'd168;
         167      :	result = 16'd168;
         168      :	result = 16'd168;
         169      :	result = 16'd169;
         170      :	result = 16'd169;
         171      :	result = 16'd169;
         172      :	result = 16'd169;
         173      :	result = 16'd169;
         174      :	result = 16'd170;
         175      :	result = 16'd170;
         176      :	result = 16'd170;
         177      :	result = 16'd170;
         178      :	result = 16'd171;
         179      :	result = 16'd171;
         180      :	result = 16'd171;
         181      :	result = 16'd171;
         182      :	result = 16'd171;
         183      :	result = 16'd172;
         184      :	result = 16'd172;
         185      :	result = 16'd172;
         186      :	result = 16'd172;
         187      :	result = 16'd172;
         188      :	result = 16'd173;
         189      :	result = 16'd173;
         190      :	result = 16'd173;
         191      :	result = 16'd173;
         192      :	result = 16'd174;
         193      :	result = 16'd174;
         194      :	result = 16'd174;
         195      :	result = 16'd174;
         196      :	result = 16'd174;
         197      :	result = 16'd175;
         198      :	result = 16'd175;
         199      :	result = 16'd175;
         200      :	result = 16'd175;
         201      :	result = 16'd176;
         202      :	result = 16'd176;
         203      :	result = 16'd176;
         204      :	result = 16'd176;
         205      :	result = 16'd176;
         206      :	result = 16'd177;
         207      :	result = 16'd177;
         208      :	result = 16'd177;
         209      :	result = 16'd177;
         210      :	result = 16'd177;
         211      :	result = 16'd178;
         212      :	result = 16'd178;
         213      :	result = 16'd178;
         214      :	result = 16'd178;
         215      :	result = 16'd179;
         216      :	result = 16'd179;
         217      :	result = 16'd179;
         218      :	result = 16'd179;
         219      :	result = 16'd179;
         220      :	result = 16'd180;
         221      :	result = 16'd180;
         222      :	result = 16'd180;
         223      :	result = 16'd180;
         224      :	result = 16'd180;
         225      :	result = 16'd181;
         226      :	result = 16'd181;
         227      :	result = 16'd181;
         228      :	result = 16'd181;
         229      :	result = 16'd181;
         230      :	result = 16'd182;
         231      :	result = 16'd182;
         232      :	result = 16'd182;
         233      :	result = 16'd182;
         234      :	result = 16'd182;
         235      :	result = 16'd183;
         236      :	result = 16'd183;
         237      :	result = 16'd183;
         238      :	result = 16'd183;
         239      :	result = 16'd183;
         240      :	result = 16'd184;
         241      :	result = 16'd184;
         242      :	result = 16'd184;
         243      :	result = 16'd184;
         244      :	result = 16'd184;
         245      :	result = 16'd185;
         246      :	result = 16'd185;
         247      :	result = 16'd185;
         248      :	result = 16'd185;
         249      :	result = 16'd185;
         250      :	result = 16'd186;
         251      :	result = 16'd186;
         252      :	result = 16'd186;
         253      :	result = 16'd186;
         254      :	result = 16'd186;
         255      :	result = 16'd187;
         256      :	result = 16'd187;
         257      :	result = 16'd187;
         258      :	result = 16'd187;
         259      :	result = 16'd187;
         260      :	result = 16'd188;
         261      :	result = 16'd188;
         262      :	result = 16'd188;
         263      :	result = 16'd188;
         264      :	result = 16'd188;
         265      :	result = 16'd189;
         266      :	result = 16'd189;
         267      :	result = 16'd189;
         268      :	result = 16'd189;
         269      :	result = 16'd189;
         270      :	result = 16'd190;
         271      :	result = 16'd190;
         272      :	result = 16'd190;
         273      :	result = 16'd190;
         274      :	result = 16'd190;
         275      :	result = 16'd191;
         276      :	result = 16'd191;
         277      :	result = 16'd191;
         278      :	result = 16'd191;
         279      :	result = 16'd191;
         280      :	result = 16'd191;
         281      :	result = 16'd192;
         282      :	result = 16'd192;
         283      :	result = 16'd192;
         284      :	result = 16'd192;
         285      :	result = 16'd192;
         286      :	result = 16'd193;
         287      :	result = 16'd193;
         288      :	result = 16'd193;
         289      :	result = 16'd193;
         290      :	result = 16'd193;
         291      :	result = 16'd193;
         292      :	result = 16'd194;
         293      :	result = 16'd194;
         294      :	result = 16'd194;
         295      :	result = 16'd194;
         296      :	result = 16'd194;
         297      :	result = 16'd195;
         298      :	result = 16'd195;
         299      :	result = 16'd195;
         300      :	result = 16'd195;
         301      :	result = 16'd195;
         302      :	result = 16'd195;
         303      :	result = 16'd196;
         304      :	result = 16'd196;
         305      :	result = 16'd196;
         306      :	result = 16'd196;
         307      :	result = 16'd196;
         308      :	result = 16'd197;
         309      :	result = 16'd197;
         310      :	result = 16'd197;
         311      :	result = 16'd197;
         312      :	result = 16'd197;
         313      :	result = 16'd197;
         314      :	result = 16'd198;
         315      :	result = 16'd198;
         316      :	result = 16'd198;
         317      :	result = 16'd198;
         318      :	result = 16'd198;
         319      :	result = 16'd198;
         320      :	result = 16'd199;
         321      :	result = 16'd199;
         322      :	result = 16'd199;
         323      :	result = 16'd199;
         324      :	result = 16'd199;
         325      :	result = 16'd200;
         326      :	result = 16'd200;
         327      :	result = 16'd200;
         328      :	result = 16'd200;
         329      :	result = 16'd200;
         330      :	result = 16'd200;
         331      :	result = 16'd201;
         332      :	result = 16'd201;
         333      :	result = 16'd201;
         334      :	result = 16'd201;
         335      :	result = 16'd201;
         336      :	result = 16'd201;
         337      :	result = 16'd202;
         338      :	result = 16'd202;
         339      :	result = 16'd202;
         340      :	result = 16'd202;
         341      :	result = 16'd202;
         342      :	result = 16'd202;
         343      :	result = 16'd203;
         344      :	result = 16'd203;
         345      :	result = 16'd203;
         346      :	result = 16'd203;
         347      :	result = 16'd203;
         348      :	result = 16'd203;
         349      :	result = 16'd204;
         350      :	result = 16'd204;
         351      :	result = 16'd204;
         352      :	result = 16'd204;
         353      :	result = 16'd204;
         354      :	result = 16'd204;
         355      :	result = 16'd204;
         356      :	result = 16'd205;
         357      :	result = 16'd205;
         358      :	result = 16'd205;
         359      :	result = 16'd205;
         360      :	result = 16'd205;
         361      :	result = 16'd205;
         362      :	result = 16'd206;
         363      :	result = 16'd206;
         364      :	result = 16'd206;
         365      :	result = 16'd206;
         366      :	result = 16'd206;
         367      :	result = 16'd206;
         368      :	result = 16'd207;
         369      :	result = 16'd207;
         370      :	result = 16'd207;
         371      :	result = 16'd207;
         372      :	result = 16'd207;
         373      :	result = 16'd207;
         374      :	result = 16'd207;
         375      :	result = 16'd208;
         376      :	result = 16'd208;
         377      :	result = 16'd208;
         378      :	result = 16'd208;
         379      :	result = 16'd208;
         380      :	result = 16'd208;
         381      :	result = 16'd209;
         382      :	result = 16'd209;
         383      :	result = 16'd209;
         384      :	result = 16'd209;
         385      :	result = 16'd209;
         386      :	result = 16'd209;
         387      :	result = 16'd209;
         388      :	result = 16'd210;
         389      :	result = 16'd210;
         390      :	result = 16'd210;
         391      :	result = 16'd210;
         392      :	result = 16'd210;
         393      :	result = 16'd210;
         394      :	result = 16'd210;
         395      :	result = 16'd211;
         396      :	result = 16'd211;
         397      :	result = 16'd211;
         398      :	result = 16'd211;
         399      :	result = 16'd211;
         400      :	result = 16'd211;
         401      :	result = 16'd211;
         402      :	result = 16'd212;
         403      :	result = 16'd212;
         404      :	result = 16'd212;
         405      :	result = 16'd212;
         406      :	result = 16'd212;
         407      :	result = 16'd212;
         408      :	result = 16'd212;
         409      :	result = 16'd213;
         410      :	result = 16'd213;
         411      :	result = 16'd213;
         412      :	result = 16'd213;
         413      :	result = 16'd213;
         414      :	result = 16'd213;
         415      :	result = 16'd213;
         416      :	result = 16'd214;
         417      :	result = 16'd214;
         418      :	result = 16'd214;
         419      :	result = 16'd214;
         420      :	result = 16'd214;
         421      :	result = 16'd214;
         422      :	result = 16'd214;
         423      :	result = 16'd214;
         424      :	result = 16'd215;
         425      :	result = 16'd215;
         426      :	result = 16'd215;
         427      :	result = 16'd215;
         428      :	result = 16'd215;
         429      :	result = 16'd215;
         430      :	result = 16'd215;
         431      :	result = 16'd216;
         432      :	result = 16'd216;
         433      :	result = 16'd216;
         434      :	result = 16'd216;
         435      :	result = 16'd216;
         436      :	result = 16'd216;
         437      :	result = 16'd216;
         438      :	result = 16'd216;
         439      :	result = 16'd217;
         440      :	result = 16'd217;
         441      :	result = 16'd217;
         442      :	result = 16'd217;
         443      :	result = 16'd217;
         444      :	result = 16'd217;
         445      :	result = 16'd217;
         446      :	result = 16'd217;
         447      :	result = 16'd218;
         448      :	result = 16'd218;
         449      :	result = 16'd218;
         450      :	result = 16'd218;
         451      :	result = 16'd218;
         452      :	result = 16'd218;
         453      :	result = 16'd218;
         454      :	result = 16'd218;
         455      :	result = 16'd219;
         456      :	result = 16'd219;
         457      :	result = 16'd219;
         458      :	result = 16'd219;
         459      :	result = 16'd219;
         460      :	result = 16'd219;
         461      :	result = 16'd219;
         462      :	result = 16'd219;
         463      :	result = 16'd220;
         464      :	result = 16'd220;
         465      :	result = 16'd220;
         466      :	result = 16'd220;
         467      :	result = 16'd220;
         468      :	result = 16'd220;
         469      :	result = 16'd220;
         470      :	result = 16'd220;
         471      :	result = 16'd221;
         472      :	result = 16'd221;
         473      :	result = 16'd221;
         474      :	result = 16'd221;
         475      :	result = 16'd221;
         476      :	result = 16'd221;
         477      :	result = 16'd221;
         478      :	result = 16'd221;
         479      :	result = 16'd221;
         480      :	result = 16'd222;
         481      :	result = 16'd222;
         482      :	result = 16'd222;
         483      :	result = 16'd222;
         484      :	result = 16'd222;
         485      :	result = 16'd222;
         486      :	result = 16'd222;
         487      :	result = 16'd222;
         488      :	result = 16'd222;
         489      :	result = 16'd223;
         490      :	result = 16'd223;
         491      :	result = 16'd223;
         492      :	result = 16'd223;
         493      :	result = 16'd223;
         494      :	result = 16'd223;
         495      :	result = 16'd223;
         496      :	result = 16'd223;
         497      :	result = 16'd223;
         498      :	result = 16'd224;
         499      :	result = 16'd224;
         500      :	result = 16'd224;
         501      :	result = 16'd224;
         502      :	result = 16'd224;
         503      :	result = 16'd224;
         504      :	result = 16'd224;
         505      :	result = 16'd224;
         506      :	result = 16'd224;
         507      :	result = 16'd225;
         508      :	result = 16'd225;
         509      :	result = 16'd225;
         510      :	result = 16'd225;
         511      :	result = 16'd225;
         512      :	result = 16'd225;
         513      :	result = 16'd225;
         514      :	result = 16'd225;
         515      :	result = 16'd225;
         516      :	result = 16'd226;
         517      :	result = 16'd226;
         518      :	result = 16'd226;
         519      :	result = 16'd226;
         520      :	result = 16'd226;
         521      :	result = 16'd226;
         522      :	result = 16'd226;
         523      :	result = 16'd226;
         524      :	result = 16'd226;
         525      :	result = 16'd226;
         526      :	result = 16'd227;
         527      :	result = 16'd227;
         528      :	result = 16'd227;
         529      :	result = 16'd227;
         530      :	result = 16'd227;
         531      :	result = 16'd227;
         532      :	result = 16'd227;
         533      :	result = 16'd227;
         534      :	result = 16'd227;
         535      :	result = 16'd227;
         536      :	result = 16'd228;
         537      :	result = 16'd228;
         538      :	result = 16'd228;
         539      :	result = 16'd228;
         540      :	result = 16'd228;
         541      :	result = 16'd228;
         542      :	result = 16'd228;
         543      :	result = 16'd228;
         544      :	result = 16'd228;
         545      :	result = 16'd228;
         546      :	result = 16'd228;
         547      :	result = 16'd229;
         548      :	result = 16'd229;
         549      :	result = 16'd229;
         550      :	result = 16'd229;
         551      :	result = 16'd229;
         552      :	result = 16'd229;
         553      :	result = 16'd229;
         554      :	result = 16'd229;
         555      :	result = 16'd229;
         556      :	result = 16'd229;
         557      :	result = 16'd229;
         558      :	result = 16'd230;
         559      :	result = 16'd230;
         560      :	result = 16'd230;
         561      :	result = 16'd230;
         562      :	result = 16'd230;
         563      :	result = 16'd230;
         564      :	result = 16'd230;
         565      :	result = 16'd230;
         566      :	result = 16'd230;
         567      :	result = 16'd230;
         568      :	result = 16'd230;
         569      :	result = 16'd231;
         570      :	result = 16'd231;
         571      :	result = 16'd231;
         572      :	result = 16'd231;
         573      :	result = 16'd231;
         574      :	result = 16'd231;
         575      :	result = 16'd231;
         576      :	result = 16'd231;
         577      :	result = 16'd231;
         578      :	result = 16'd231;
         579      :	result = 16'd231;
         580      :	result = 16'd232;
         581      :	result = 16'd232;
         582      :	result = 16'd232;
         583      :	result = 16'd232;
         584      :	result = 16'd232;
         585      :	result = 16'd232;
         586      :	result = 16'd232;
         587      :	result = 16'd232;
         588      :	result = 16'd232;
         589      :	result = 16'd232;
         590      :	result = 16'd232;
         591      :	result = 16'd232;
         592      :	result = 16'd233;
         593      :	result = 16'd233;
         594      :	result = 16'd233;
         595      :	result = 16'd233;
         596      :	result = 16'd233;
         597      :	result = 16'd233;
         598      :	result = 16'd233;
         599      :	result = 16'd233;
         600      :	result = 16'd233;
         601      :	result = 16'd233;
         602      :	result = 16'd233;
         603      :	result = 16'd233;
         604      :	result = 16'd233;
         605      :	result = 16'd234;
         606      :	result = 16'd234;
         607      :	result = 16'd234;
         608      :	result = 16'd234;
         609      :	result = 16'd234;
         610      :	result = 16'd234;
         611      :	result = 16'd234;
         612      :	result = 16'd234;
         613      :	result = 16'd234;
         614      :	result = 16'd234;
         615      :	result = 16'd234;
         616      :	result = 16'd234;
         617      :	result = 16'd234;
         618      :	result = 16'd235;
         619      :	result = 16'd235;
         620      :	result = 16'd235;
         621      :	result = 16'd235;
         622      :	result = 16'd235;
         623      :	result = 16'd235;
         624      :	result = 16'd235;
         625      :	result = 16'd235;
         626      :	result = 16'd235;
         627      :	result = 16'd235;
         628      :	result = 16'd235;
         629      :	result = 16'd235;
         630      :	result = 16'd235;
         631      :	result = 16'd236;
         632      :	result = 16'd236;
         633      :	result = 16'd236;
         634      :	result = 16'd236;
         635      :	result = 16'd236;
         636      :	result = 16'd236;
         637      :	result = 16'd236;
         638      :	result = 16'd236;
         639      :	result = 16'd236;
         640      :	result = 16'd236;
         641      :	result = 16'd236;
         642      :	result = 16'd236;
         643      :	result = 16'd236;
         644      :	result = 16'd236;
         645      :	result = 16'd236;
         646      :	result = 16'd237;
         647      :	result = 16'd237;
         648      :	result = 16'd237;
         649      :	result = 16'd237;
         650      :	result = 16'd237;
         651      :	result = 16'd237;
         652      :	result = 16'd237;
         653      :	result = 16'd237;
         654      :	result = 16'd237;
         655      :	result = 16'd237;
         656      :	result = 16'd237;
         657      :	result = 16'd237;
         658      :	result = 16'd237;
         659      :	result = 16'd237;
         660      :	result = 16'd238;
         661      :	result = 16'd238;
         662      :	result = 16'd238;
         663      :	result = 16'd238;
         664      :	result = 16'd238;
         665      :	result = 16'd238;
         666      :	result = 16'd238;
         667      :	result = 16'd238;
         668      :	result = 16'd238;
         669      :	result = 16'd238;
         670      :	result = 16'd238;
         671      :	result = 16'd238;
         672      :	result = 16'd238;
         673      :	result = 16'd238;
         674      :	result = 16'd238;
         675      :	result = 16'd238;
         676      :	result = 16'd239;
         677      :	result = 16'd239;
         678      :	result = 16'd239;
         679      :	result = 16'd239;
         680      :	result = 16'd239;
         681      :	result = 16'd239;
         682      :	result = 16'd239;
         683      :	result = 16'd239;
         684      :	result = 16'd239;
         685      :	result = 16'd239;
         686      :	result = 16'd239;
         687      :	result = 16'd239;
         688      :	result = 16'd239;
         689      :	result = 16'd239;
         690      :	result = 16'd239;
         691      :	result = 16'd239;
         692      :	result = 16'd239;
         693      :	result = 16'd240;
         694      :	result = 16'd240;
         695      :	result = 16'd240;
         696      :	result = 16'd240;
         697      :	result = 16'd240;
         698      :	result = 16'd240;
         699      :	result = 16'd240;
         700      :	result = 16'd240;
         701      :	result = 16'd240;
         702      :	result = 16'd240;
         703      :	result = 16'd240;
         704      :	result = 16'd240;
         705      :	result = 16'd240;
         706      :	result = 16'd240;
         707      :	result = 16'd240;
         708      :	result = 16'd240;
         709      :	result = 16'd240;
         710      :	result = 16'd241;
         711      :	result = 16'd241;
         712      :	result = 16'd241;
         713      :	result = 16'd241;
         714      :	result = 16'd241;
         715      :	result = 16'd241;
         716      :	result = 16'd241;
         717      :	result = 16'd241;
         718      :	result = 16'd241;
         719      :	result = 16'd241;
         720      :	result = 16'd241;
         721      :	result = 16'd241;
         722      :	result = 16'd241;
         723      :	result = 16'd241;
         724      :	result = 16'd241;
         725      :	result = 16'd241;
         726      :	result = 16'd241;
         727      :	result = 16'd241;
         728      :	result = 16'd241;
         729      :	result = 16'd242;
         730      :	result = 16'd242;
         731      :	result = 16'd242;
         732      :	result = 16'd242;
         733      :	result = 16'd242;
         734      :	result = 16'd242;
         735      :	result = 16'd242;
         736      :	result = 16'd242;
         737      :	result = 16'd242;
         738      :	result = 16'd242;
         739      :	result = 16'd242;
         740      :	result = 16'd242;
         741      :	result = 16'd242;
         742      :	result = 16'd242;
         743      :	result = 16'd242;
         744      :	result = 16'd242;
         745      :	result = 16'd242;
         746      :	result = 16'd242;
         747      :	result = 16'd242;
         748      :	result = 16'd242;
         749      :	result = 16'd243;
         750      :	result = 16'd243;
         751      :	result = 16'd243;
         752      :	result = 16'd243;
         753      :	result = 16'd243;
         754      :	result = 16'd243;
         755      :	result = 16'd243;
         756      :	result = 16'd243;
         757      :	result = 16'd243;
         758      :	result = 16'd243;
         759      :	result = 16'd243;
         760      :	result = 16'd243;
         761      :	result = 16'd243;
         762      :	result = 16'd243;
         763      :	result = 16'd243;
         764      :	result = 16'd243;
         765      :	result = 16'd243;
         766      :	result = 16'd243;
         767      :	result = 16'd243;
         768      :	result = 16'd243;
         769      :	result = 16'd243;
         770      :	result = 16'd243;
         771      :	result = 16'd244;
         772      :	result = 16'd244;
         773      :	result = 16'd244;
         774      :	result = 16'd244;
         775      :	result = 16'd244;
         776      :	result = 16'd244;
         777      :	result = 16'd244;
         778      :	result = 16'd244;
         779      :	result = 16'd244;
         780      :	result = 16'd244;
         781      :	result = 16'd244;
         782      :	result = 16'd244;
         783      :	result = 16'd244;
         784      :	result = 16'd244;
         785      :	result = 16'd244;
         786      :	result = 16'd244;
         787      :	result = 16'd244;
         788      :	result = 16'd244;
         789      :	result = 16'd244;
         790      :	result = 16'd244;
         791      :	result = 16'd244;
         792      :	result = 16'd244;
         793      :	result = 16'd244;
         794      :	result = 16'd245;
         795      :	result = 16'd245;
         796      :	result = 16'd245;
         797      :	result = 16'd245;
         798      :	result = 16'd245;
         799      :	result = 16'd245;
         800      :	result = 16'd245;
         801      :	result = 16'd245;
         802      :	result = 16'd245;
         803      :	result = 16'd245;
         804      :	result = 16'd245;
         805      :	result = 16'd245;
         806      :	result = 16'd245;
         807      :	result = 16'd245;
         808      :	result = 16'd245;
         809      :	result = 16'd245;
         810      :	result = 16'd245;
         811      :	result = 16'd245;
         812      :	result = 16'd245;
         813      :	result = 16'd245;
         814      :	result = 16'd245;
         815      :	result = 16'd245;
         816      :	result = 16'd245;
         817      :	result = 16'd245;
         818      :	result = 16'd245;
         819      :	result = 16'd246;
         820      :	result = 16'd246;
         821      :	result = 16'd246;
         822      :	result = 16'd246;
         823      :	result = 16'd246;
         824      :	result = 16'd246;
         825      :	result = 16'd246;
         826      :	result = 16'd246;
         827      :	result = 16'd246;
         828      :	result = 16'd246;
         829      :	result = 16'd246;
         830      :	result = 16'd246;
         831      :	result = 16'd246;
         832      :	result = 16'd246;
         833      :	result = 16'd246;
         834      :	result = 16'd246;
         835      :	result = 16'd246;
         836      :	result = 16'd246;
         837      :	result = 16'd246;
         838      :	result = 16'd246;
         839      :	result = 16'd246;
         840      :	result = 16'd246;
         841      :	result = 16'd246;
         842      :	result = 16'd246;
         843      :	result = 16'd246;
         844      :	result = 16'd246;
         845      :	result = 16'd246;
         846      :	result = 16'd246;
         847      :	result = 16'd247;
         848      :	result = 16'd247;
         849      :	result = 16'd247;
         850      :	result = 16'd247;
         851      :	result = 16'd247;
         852      :	result = 16'd247;
         853      :	result = 16'd247;
         854      :	result = 16'd247;
         855      :	result = 16'd247;
         856      :	result = 16'd247;
         857      :	result = 16'd247;
         858      :	result = 16'd247;
         859      :	result = 16'd247;
         860      :	result = 16'd247;
         861      :	result = 16'd247;
         862      :	result = 16'd247;
         863      :	result = 16'd247;
         864      :	result = 16'd247;
         865      :	result = 16'd247;
         866      :	result = 16'd247;
         867      :	result = 16'd247;
         868      :	result = 16'd247;
         869      :	result = 16'd247;
         870      :	result = 16'd247;
         871      :	result = 16'd247;
         872      :	result = 16'd247;
         873      :	result = 16'd247;
         874      :	result = 16'd247;
         875      :	result = 16'd247;
         876      :	result = 16'd247;
         877      :	result = 16'd247;
         878      :	result = 16'd247;
         879      :	result = 16'd248;
         880      :	result = 16'd248;
         881      :	result = 16'd248;
         882      :	result = 16'd248;
         883      :	result = 16'd248;
         884      :	result = 16'd248;
         885      :	result = 16'd248;
         886      :	result = 16'd248;
         887      :	result = 16'd248;
         888      :	result = 16'd248;
         889      :	result = 16'd248;
         890      :	result = 16'd248;
         891      :	result = 16'd248;
         892      :	result = 16'd248;
         893      :	result = 16'd248;
         894      :	result = 16'd248;
         895      :	result = 16'd248;
         896      :	result = 16'd248;
         897      :	result = 16'd248;
         898      :	result = 16'd248;
         899      :	result = 16'd248;
         900      :	result = 16'd248;
         901      :	result = 16'd248;
         902      :	result = 16'd248;
         903      :	result = 16'd248;
         904      :	result = 16'd248;
         905      :	result = 16'd248;
         906      :	result = 16'd248;
         907      :	result = 16'd248;
         908      :	result = 16'd248;
         909      :	result = 16'd248;
         910      :	result = 16'd248;
         911      :	result = 16'd248;
         912      :	result = 16'd248;
         913      :	result = 16'd248;
         914      :	result = 16'd249;
         915      :	result = 16'd249;
         916      :	result = 16'd249;
         917      :	result = 16'd249;
         918      :	result = 16'd249;
         919      :	result = 16'd249;
         920      :	result = 16'd249;
         921      :	result = 16'd249;
         922      :	result = 16'd249;
         923      :	result = 16'd249;
         924      :	result = 16'd249;
         925      :	result = 16'd249;
         926      :	result = 16'd249;
         927      :	result = 16'd249;
         928      :	result = 16'd249;
         929      :	result = 16'd249;
         930      :	result = 16'd249;
         931      :	result = 16'd249;
         932      :	result = 16'd249;
         933      :	result = 16'd249;
         934      :	result = 16'd249;
         935      :	result = 16'd249;
         936      :	result = 16'd249;
         937      :	result = 16'd249;
         938      :	result = 16'd249;
         939      :	result = 16'd249;
         940      :	result = 16'd249;
         941      :	result = 16'd249;
         942      :	result = 16'd249;
         943      :	result = 16'd249;
         944      :	result = 16'd249;
         945      :	result = 16'd249;
         946      :	result = 16'd249;
         947      :	result = 16'd249;
         948      :	result = 16'd249;
         949      :	result = 16'd249;
         950      :	result = 16'd249;
         951      :	result = 16'd249;
         952      :	result = 16'd249;
         953      :	result = 16'd249;
         954      :	result = 16'd250;
         955      :	result = 16'd250;
         956      :	result = 16'd250;
         957      :	result = 16'd250;
         958      :	result = 16'd250;
         959      :	result = 16'd250;
         960      :	result = 16'd250;
         961      :	result = 16'd250;
         962      :	result = 16'd250;
         963      :	result = 16'd250;
         964      :	result = 16'd250;
         965      :	result = 16'd250;
         966      :	result = 16'd250;
         967      :	result = 16'd250;
         968      :	result = 16'd250;
         969      :	result = 16'd250;
         970      :	result = 16'd250;
         971      :	result = 16'd250;
         972      :	result = 16'd250;
         973      :	result = 16'd250;
         974      :	result = 16'd250;
         975      :	result = 16'd250;
         976      :	result = 16'd250;
         977      :	result = 16'd250;
         978      :	result = 16'd250;
         979      :	result = 16'd250;
         980      :	result = 16'd250;
         981      :	result = 16'd250;
         982      :	result = 16'd250;
         983      :	result = 16'd250;
         984      :	result = 16'd250;
         985      :	result = 16'd250;
         986      :	result = 16'd250;
         987      :	result = 16'd250;
         988      :	result = 16'd250;
         989      :	result = 16'd250;
         990      :	result = 16'd250;
         991      :	result = 16'd250;
         992      :	result = 16'd250;
         993      :	result = 16'd250;
         994      :	result = 16'd250;
         995      :	result = 16'd250;
         996      :	result = 16'd250;
         997      :	result = 16'd250;
         998      :	result = 16'd250;
         999      :	result = 16'd250;
         1000     :	result = 16'd250;
         1001     :	result = 16'd250;
         1002     :	result = 16'd251;
         1003     :	result = 16'd251;
         1004     :	result = 16'd251;
         1005     :	result = 16'd251;
         1006     :	result = 16'd251;
         1007     :	result = 16'd251;
         1008     :	result = 16'd251;
         1009     :	result = 16'd251;
         1010     :	result = 16'd251;
         1011     :	result = 16'd251;
         1012     :	result = 16'd251;
         1013     :	result = 16'd251;
         1014     :	result = 16'd251;
         1015     :	result = 16'd251;
         1016     :	result = 16'd251;
         1017     :	result = 16'd251;
         1018     :	result = 16'd251;
         1019     :	result = 16'd251;
         1020     :	result = 16'd251;
         1021     :	result = 16'd251;
         1022     :	result = 16'd251;
         1023     :	result = 16'd251;
         1024     :	result = 16'd251;
         1025     :	result = 16'd251;
         1026     :	result = 16'd251;
         1027     :	result = 16'd251;
         1028     :	result = 16'd251;
         1029     :	result = 16'd251;
         1030     :	result = 16'd251;
         1031     :	result = 16'd251;
         1032     :	result = 16'd251;
         1033     :	result = 16'd251;
         1034     :	result = 16'd251;
         1035     :	result = 16'd251;
         1036     :	result = 16'd251;
         1037     :	result = 16'd251;
         1038     :	result = 16'd251;
         1039     :	result = 16'd251;
         1040     :	result = 16'd251;
         1041     :	result = 16'd251;
         1042     :	result = 16'd251;
         1043     :	result = 16'd251;
         1044     :	result = 16'd251;
         1045     :	result = 16'd251;
         1046     :	result = 16'd251;
         1047     :	result = 16'd251;
         1048     :	result = 16'd251;
         1049     :	result = 16'd251;
         1050     :	result = 16'd251;
         1051     :	result = 16'd251;
         1052     :	result = 16'd251;
         1053     :	result = 16'd251;
         1054     :	result = 16'd251;
         1055     :	result = 16'd251;
         1056     :	result = 16'd251;
         1057     :	result = 16'd251;
         1058     :	result = 16'd251;
         1059     :	result = 16'd251;
         1060     :	result = 16'd252;
         1061     :	result = 16'd252;
         1062     :	result = 16'd252;
         1063     :	result = 16'd252;
         1064     :	result = 16'd252;
         1065     :	result = 16'd252;
         1066     :	result = 16'd252;
         1067     :	result = 16'd252;
         1068     :	result = 16'd252;
         1069     :	result = 16'd252;
         1070     :	result = 16'd252;
         1071     :	result = 16'd252;
         1072     :	result = 16'd252;
         1073     :	result = 16'd252;
         1074     :	result = 16'd252;
         1075     :	result = 16'd252;
         1076     :	result = 16'd252;
         1077     :	result = 16'd252;
         1078     :	result = 16'd252;
         1079     :	result = 16'd252;
         1080     :	result = 16'd252;
         1081     :	result = 16'd252;
         1082     :	result = 16'd252;
         1083     :	result = 16'd252;
         1084     :	result = 16'd252;
         1085     :	result = 16'd252;
         1086     :	result = 16'd252;
         1087     :	result = 16'd252;
         1088     :	result = 16'd252;
         1089     :	result = 16'd252;
         1090     :	result = 16'd252;
         1091     :	result = 16'd252;
         1092     :	result = 16'd252;
         1093     :	result = 16'd252;
         1094     :	result = 16'd252;
         1095     :	result = 16'd252;
         1096     :	result = 16'd252;
         1097     :	result = 16'd252;
         1098     :	result = 16'd252;
         1099     :	result = 16'd252;
         1100     :	result = 16'd252;
         1101     :	result = 16'd252;
         1102     :	result = 16'd252;
         1103     :	result = 16'd252;
         1104     :	result = 16'd252;
         1105     :	result = 16'd252;
         1106     :	result = 16'd252;
         1107     :	result = 16'd252;
         1108     :	result = 16'd252;
         1109     :	result = 16'd252;
         1110     :	result = 16'd252;
         1111     :	result = 16'd252;
         1112     :	result = 16'd252;
         1113     :	result = 16'd252;
         1114     :	result = 16'd252;
         1115     :	result = 16'd252;
         1116     :	result = 16'd252;
         1117     :	result = 16'd252;
         1118     :	result = 16'd252;
         1119     :	result = 16'd252;
         1120     :	result = 16'd252;
         1121     :	result = 16'd252;
         1122     :	result = 16'd252;
         1123     :	result = 16'd252;
         1124     :	result = 16'd252;
         1125     :	result = 16'd252;
         1126     :	result = 16'd252;
         1127     :	result = 16'd252;
         1128     :	result = 16'd252;
         1129     :	result = 16'd252;
         1130     :	result = 16'd252;
         1131     :	result = 16'd252;
         1132     :	result = 16'd252;
         1133     :	result = 16'd252;
         1134     :	result = 16'd252;
         1135     :	result = 16'd253;
         1136     :	result = 16'd253;
         1137     :	result = 16'd253;
         1138     :	result = 16'd253;
         1139     :	result = 16'd253;
         1140     :	result = 16'd253;
         1141     :	result = 16'd253;
         1142     :	result = 16'd253;
         1143     :	result = 16'd253;
         1144     :	result = 16'd253;
         1145     :	result = 16'd253;
         1146     :	result = 16'd253;
         1147     :	result = 16'd253;
         1148     :	result = 16'd253;
         1149     :	result = 16'd253;
         1150     :	result = 16'd253;
         1151     :	result = 16'd253;
         1152     :	result = 16'd253;
         1153     :	result = 16'd253;
         1154     :	result = 16'd253;
         1155     :	result = 16'd253;
         1156     :	result = 16'd253;
         1157     :	result = 16'd253;
         1158     :	result = 16'd253;
         1159     :	result = 16'd253;
         1160     :	result = 16'd253;
         1161     :	result = 16'd253;
         1162     :	result = 16'd253;
         1163     :	result = 16'd253;
         1164     :	result = 16'd253;
         1165     :	result = 16'd253;
         1166     :	result = 16'd253;
         1167     :	result = 16'd253;
         1168     :	result = 16'd253;
         1169     :	result = 16'd253;
         1170     :	result = 16'd253;
         1171     :	result = 16'd253;
         1172     :	result = 16'd253;
         1173     :	result = 16'd253;
         1174     :	result = 16'd253;
         1175     :	result = 16'd253;
         1176     :	result = 16'd253;
         1177     :	result = 16'd253;
         1178     :	result = 16'd253;
         1179     :	result = 16'd253;
         1180     :	result = 16'd253;
         1181     :	result = 16'd253;
         1182     :	result = 16'd253;
         1183     :	result = 16'd253;
         1184     :	result = 16'd253;
         1185     :	result = 16'd253;
         1186     :	result = 16'd253;
         1187     :	result = 16'd253;
         1188     :	result = 16'd253;
         1189     :	result = 16'd253;
         1190     :	result = 16'd253;
         1191     :	result = 16'd253;
         1192     :	result = 16'd253;
         1193     :	result = 16'd253;
         1194     :	result = 16'd253;
         1195     :	result = 16'd253;
         1196     :	result = 16'd253;
         1197     :	result = 16'd253;
         1198     :	result = 16'd253;
         1199     :	result = 16'd253;
         1200     :	result = 16'd253;
         1201     :	result = 16'd253;
         1202     :	result = 16'd253;
         1203     :	result = 16'd253;
         1204     :	result = 16'd253;
         1205     :	result = 16'd253;
         1206     :	result = 16'd253;
         1207     :	result = 16'd253;
         1208     :	result = 16'd253;
         1209     :	result = 16'd253;
         1210     :	result = 16'd253;
         1211     :	result = 16'd253;
         1212     :	result = 16'd253;
         1213     :	result = 16'd253;
         1214     :	result = 16'd253;
         1215     :	result = 16'd253;
         1216     :	result = 16'd253;
         1217     :	result = 16'd253;
         1218     :	result = 16'd253;
         1219     :	result = 16'd253;
         1220     :	result = 16'd253;
         1221     :	result = 16'd253;
         1222     :	result = 16'd253;
         1223     :	result = 16'd253;
         1224     :	result = 16'd253;
         1225     :	result = 16'd253;
         1226     :	result = 16'd253;
         1227     :	result = 16'd253;
         1228     :	result = 16'd253;
         1229     :	result = 16'd253;
         1230     :	result = 16'd253;
         1231     :	result = 16'd253;
         1232     :	result = 16'd253;
         1233     :	result = 16'd253;
         1234     :	result = 16'd253;
         1235     :	result = 16'd253;
         1236     :	result = 16'd253;
         1237     :	result = 16'd253;
         1238     :	result = 16'd253;
         1239     :	result = 16'd253;
         1240     :	result = 16'd254;
         1241     :	result = 16'd254;
         1242     :	result = 16'd254;
         1243     :	result = 16'd254;
         1244     :	result = 16'd254;
         1245     :	result = 16'd254;
         1246     :	result = 16'd254;
         1247     :	result = 16'd254;
         1248     :	result = 16'd254;
         1249     :	result = 16'd254;
         1250     :	result = 16'd254;
         1251     :	result = 16'd254;
         1252     :	result = 16'd254;
         1253     :	result = 16'd254;
         1254     :	result = 16'd254;
         1255     :	result = 16'd254;
         1256     :	result = 16'd254;
         1257     :	result = 16'd254;
         1258     :	result = 16'd254;
         1259     :	result = 16'd254;
         1260     :	result = 16'd254;
         1261     :	result = 16'd254;
         1262     :	result = 16'd254;
         1263     :	result = 16'd254;
         1264     :	result = 16'd254;
         1265     :	result = 16'd254;
         1266     :	result = 16'd254;
         1267     :	result = 16'd254;
         1268     :	result = 16'd254;
         1269     :	result = 16'd254;
         1270     :	result = 16'd254;
         1271     :	result = 16'd254;
         1272     :	result = 16'd254;
         1273     :	result = 16'd254;
         1274     :	result = 16'd254;
         1275     :	result = 16'd254;
         1276     :	result = 16'd254;
         1277     :	result = 16'd254;
         1278     :	result = 16'd254;
         1279     :	result = 16'd254;
         1280     :	result = 16'd254;
         1281     :	result = 16'd254;
         1282     :	result = 16'd254;
         1283     :	result = 16'd254;
         1284     :	result = 16'd254;
         1285     :	result = 16'd254;
         1286     :	result = 16'd254;
         1287     :	result = 16'd254;
         1288     :	result = 16'd254;
         1289     :	result = 16'd254;
         1290     :	result = 16'd254;
         1291     :	result = 16'd254;
         1292     :	result = 16'd254;
         1293     :	result = 16'd254;
         1294     :	result = 16'd254;
         1295     :	result = 16'd254;
         1296     :	result = 16'd254;
         1297     :	result = 16'd254;
         1298     :	result = 16'd254;
         1299     :	result = 16'd254;
         1300     :	result = 16'd254;
         1301     :	result = 16'd254;
         1302     :	result = 16'd254;
         1303     :	result = 16'd254;
         1304     :	result = 16'd254;
         1305     :	result = 16'd254;
         1306     :	result = 16'd254;
         1307     :	result = 16'd254;
         1308     :	result = 16'd254;
         1309     :	result = 16'd254;
         1310     :	result = 16'd254;
         1311     :	result = 16'd254;
         1312     :	result = 16'd254;
         1313     :	result = 16'd254;
         1314     :	result = 16'd254;
         1315     :	result = 16'd254;
         1316     :	result = 16'd254;
         1317     :	result = 16'd254;
         1318     :	result = 16'd254;
         1319     :	result = 16'd254;
         1320     :	result = 16'd254;
         1321     :	result = 16'd254;
         1322     :	result = 16'd254;
         1323     :	result = 16'd254;
         1324     :	result = 16'd254;
         1325     :	result = 16'd254;
         1326     :	result = 16'd254;
         1327     :	result = 16'd254;
         1328     :	result = 16'd254;
         1329     :	result = 16'd254;
         1330     :	result = 16'd254;
         1331     :	result = 16'd254;
         1332     :	result = 16'd254;
         1333     :	result = 16'd254;
         1334     :	result = 16'd254;
         1335     :	result = 16'd254;
         1336     :	result = 16'd254;
         1337     :	result = 16'd254;
         1338     :	result = 16'd254;
         1339     :	result = 16'd254;
         1340     :	result = 16'd254;
         1341     :	result = 16'd254;
         1342     :	result = 16'd254;
         1343     :	result = 16'd254;
         1344     :	result = 16'd254;
         1345     :	result = 16'd254;
         1346     :	result = 16'd254;
         1347     :	result = 16'd254;
         1348     :	result = 16'd254;
         1349     :	result = 16'd254;
         1350     :	result = 16'd254;
         1351     :	result = 16'd254;
         1352     :	result = 16'd254;
         1353     :	result = 16'd254;
         1354     :	result = 16'd254;
         1355     :	result = 16'd254;
         1356     :	result = 16'd254;
         1357     :	result = 16'd254;
         1358     :	result = 16'd254;
         1359     :	result = 16'd254;
         1360     :	result = 16'd254;
         1361     :	result = 16'd254;
         1362     :	result = 16'd254;
         1363     :	result = 16'd254;
         1364     :	result = 16'd254;
         1365     :	result = 16'd254;
         1366     :	result = 16'd254;
         1367     :	result = 16'd254;
         1368     :	result = 16'd254;
         1369     :	result = 16'd254;
         1370     :	result = 16'd254;
         1371     :	result = 16'd254;
         1372     :	result = 16'd254;
         1373     :	result = 16'd254;
         1374     :	result = 16'd254;
         1375     :	result = 16'd254;
         1376     :	result = 16'd254;
         1377     :	result = 16'd254;
         1378     :	result = 16'd254;
         1379     :	result = 16'd254;
         1380     :	result = 16'd254;
         1381     :	result = 16'd254;
         1382     :	result = 16'd254;
         1383     :	result = 16'd254;
         1384     :	result = 16'd254;
         1385     :	result = 16'd254;
         1386     :	result = 16'd254;
         1387     :	result = 16'd254;
         1388     :	result = 16'd254;
         1389     :	result = 16'd254;
         1390     :	result = 16'd254;
         1391     :	result = 16'd254;
         1392     :	result = 16'd254;
         1393     :	result = 16'd254;
         1394     :	result = 16'd254;
         1395     :	result = 16'd254;
         1396     :	result = 16'd254;
         1397     :	result = 16'd254;
         1398     :	result = 16'd254;
         1399     :	result = 16'd254;
         1400     :	result = 16'd254;
         1401     :	result = 16'd254;
         1402     :	result = 16'd254;
         1403     :	result = 16'd254;
         1404     :	result = 16'd254;
         1405     :	result = 16'd254;
         1406     :	result = 16'd254;
         1407     :	result = 16'd254;
         1408     :	result = 16'd254;
         1409     :	result = 16'd254;
         1410     :	result = 16'd254;
         1411     :	result = 16'd254;
         1412     :	result = 16'd254;
         1413     :	result = 16'd254;
         1414     :	result = 16'd254;
         1415     :	result = 16'd254;
         1416     :	result = 16'd254;
         1417     :	result = 16'd254;
         1418     :	result = 16'd255;
         1419     :	result = 16'd255;
         1420     :	result = 16'd255;
         1421     :	result = 16'd255;
         1422     :	result = 16'd255;
         1423     :	result = 16'd255;
         1424     :	result = 16'd255;
         1425     :	result = 16'd255;
         1426     :	result = 16'd255;
         1427     :	result = 16'd255;
         1428     :	result = 16'd255;
         1429     :	result = 16'd255;
         1430     :	result = 16'd255;
         1431     :	result = 16'd255;
         1432     :	result = 16'd255;
         1433     :	result = 16'd255;
         1434     :	result = 16'd255;
         1435     :	result = 16'd255;
         1436     :	result = 16'd255;
         1437     :	result = 16'd255;
         1438     :	result = 16'd255;
         1439     :	result = 16'd255;
         1440     :	result = 16'd255;
         1441     :	result = 16'd255;
         1442     :	result = 16'd255;
         1443     :	result = 16'd255;
         1444     :	result = 16'd255;
         1445     :	result = 16'd255;
         1446     :	result = 16'd255;
         1447     :	result = 16'd255;
         1448     :	result = 16'd255;
         1449     :	result = 16'd255;
         1450     :	result = 16'd255;
         1451     :	result = 16'd255;
         1452     :	result = 16'd255;
         1453     :	result = 16'd255;
         1454     :	result = 16'd255;
         1455     :	result = 16'd255;
         1456     :	result = 16'd255;
         1457     :	result = 16'd255;
         1458     :	result = 16'd255;
         1459     :	result = 16'd255;
         1460     :	result = 16'd255;
         1461     :	result = 16'd255;
         1462     :	result = 16'd255;
         1463     :	result = 16'd255;
         1464     :	result = 16'd255;
         1465     :	result = 16'd255;
         1466     :	result = 16'd255;
         1467     :	result = 16'd255;
         1468     :	result = 16'd255;
         1469     :	result = 16'd255;
         1470     :	result = 16'd255;
         1471     :	result = 16'd255;
         1472     :	result = 16'd255;
         1473     :	result = 16'd255;
         1474     :	result = 16'd255;
         1475     :	result = 16'd255;
         1476     :	result = 16'd255;
         1477     :	result = 16'd255;
         1478     :	result = 16'd255;
         1479     :	result = 16'd255;
         1480     :	result = 16'd255;
         1481     :	result = 16'd255;
         1482     :	result = 16'd255;
         1483     :	result = 16'd255;
         1484     :	result = 16'd255;
         1485     :	result = 16'd255;
         1486     :	result = 16'd255;
         1487     :	result = 16'd255;
         1488     :	result = 16'd255;
         1489     :	result = 16'd255;
         1490     :	result = 16'd255;
         1491     :	result = 16'd255;
         1492     :	result = 16'd255;
         1493     :	result = 16'd255;
         1494     :	result = 16'd255;
         1495     :	result = 16'd255;
         1496     :	result = 16'd255;
         1497     :	result = 16'd255;
         1498     :	result = 16'd255;
         1499     :	result = 16'd255;
         1500     :	result = 16'd255;
         1501     :	result = 16'd255;
         1502     :	result = 16'd255;
         1503     :	result = 16'd255;
         1504     :	result = 16'd255;
         1505     :	result = 16'd255;
         1506     :	result = 16'd255;
         1507     :	result = 16'd255;
         1508     :	result = 16'd255;
         1509     :	result = 16'd255;
         1510     :	result = 16'd255;
         1511     :	result = 16'd255;
         1512     :	result = 16'd255;
         1513     :	result = 16'd255;
         1514     :	result = 16'd255;
         1515     :	result = 16'd255;
         1516     :	result = 16'd255;
         1517     :	result = 16'd255;
         1518     :	result = 16'd255;
         1519     :	result = 16'd255;
         1520     :	result = 16'd255;
         1521     :	result = 16'd255;
         1522     :	result = 16'd255;
         1523     :	result = 16'd255;
         1524     :	result = 16'd255;
         1525     :	result = 16'd255;
         1526     :	result = 16'd255;
         1527     :	result = 16'd255;
         1528     :	result = 16'd255;
         1529     :	result = 16'd255;
         1530     :	result = 16'd255;
         1531     :	result = 16'd255;
         1532     :	result = 16'd255;
         1533     :	result = 16'd255;
         1534     :	result = 16'd255;
         1535     :	result = 16'd255;
         1536     :	result = 16'd255;
         1537     :	result = 16'd255;
         1538     :	result = 16'd255;
         1539     :	result = 16'd255;
         1540     :	result = 16'd255;
         1541     :	result = 16'd255;
         1542     :	result = 16'd255;
         1543     :	result = 16'd255;
         1544     :	result = 16'd255;
         1545     :	result = 16'd255;
         1546     :	result = 16'd255;
         1547     :	result = 16'd255;
         1548     :	result = 16'd255;
         1549     :	result = 16'd255;
         1550     :	result = 16'd255;
         1551     :	result = 16'd255;
         1552     :	result = 16'd255;
         1553     :	result = 16'd255;
         1554     :	result = 16'd255;
         1555     :	result = 16'd255;
         1556     :	result = 16'd255;
         1557     :	result = 16'd255;
         1558     :	result = 16'd255;
         1559     :	result = 16'd255;
         1560     :	result = 16'd255;
         1561     :	result = 16'd255;
         1562     :	result = 16'd255;
         1563     :	result = 16'd255;
         1564     :	result = 16'd255;
         1565     :	result = 16'd255;
         1566     :	result = 16'd255;
         1567     :	result = 16'd255;
         1568     :	result = 16'd255;
         1569     :	result = 16'd255;
         1570     :	result = 16'd255;
         1571     :	result = 16'd255;
         1572     :	result = 16'd255;
         1573     :	result = 16'd255;
         1574     :	result = 16'd255;
         1575     :	result = 16'd255;
         1576     :	result = 16'd255;
         1577     :	result = 16'd255;
         1578     :	result = 16'd255;
         1579     :	result = 16'd255;
         1580     :	result = 16'd255;
         1581     :	result = 16'd255;
         1582     :	result = 16'd255;
         1583     :	result = 16'd255;
         1584     :	result = 16'd255;
         1585     :	result = 16'd255;
         1586     :	result = 16'd255;
         1587     :	result = 16'd255;
         1588     :	result = 16'd255;
         1589     :	result = 16'd255;
         1590     :	result = 16'd255;
         1591     :	result = 16'd255;
         1592     :	result = 16'd255;
         1593     :	result = 16'd255;
         1594     :	result = 16'd255;
         1595     :	result = 16'd255;
         1596     :	result = 16'd255;
         1597     :	result = 16'd255;
         1598     :	result = 16'd255;
         1599     :	result = 16'd255;
         1600     :	result = 16'd255;
         1601     :	result = 16'd255;
         1602     :	result = 16'd255;
         1603     :	result = 16'd255;
         1604     :	result = 16'd255;
         1605     :	result = 16'd255;
         1606     :	result = 16'd255;
         1607     :	result = 16'd255;
         1608     :	result = 16'd255;
         1609     :	result = 16'd255;
         1610     :	result = 16'd255;
         1611     :	result = 16'd255;
         1612     :	result = 16'd255;
         1613     :	result = 16'd255;
         1614     :	result = 16'd255;
         1615     :	result = 16'd255;
         1616     :	result = 16'd255;
         1617     :	result = 16'd255;
         1618     :	result = 16'd255;
         1619     :	result = 16'd255;
         1620     :	result = 16'd255;
         1621     :	result = 16'd255;
         1622     :	result = 16'd255;
         1623     :	result = 16'd255;
         1624     :	result = 16'd255;
         1625     :	result = 16'd255;
         1626     :	result = 16'd255;
         1627     :	result = 16'd255;
         1628     :	result = 16'd255;
         1629     :	result = 16'd255;
         1630     :	result = 16'd255;
         1631     :	result = 16'd255;
         1632     :	result = 16'd255;
         1633     :	result = 16'd255;
         1634     :	result = 16'd255;
         1635     :	result = 16'd255;
         1636     :	result = 16'd255;
         1637     :	result = 16'd255;
         1638     :	result = 16'd255;
         1639     :	result = 16'd255;
         1640     :	result = 16'd255;
         1641     :	result = 16'd255;
         1642     :	result = 16'd255;
         1643     :	result = 16'd255;
         1644     :	result = 16'd255;
         1645     :	result = 16'd255;
         1646     :	result = 16'd255;
         1647     :	result = 16'd255;
         1648     :	result = 16'd255;
         1649     :	result = 16'd255;
         1650     :	result = 16'd255;
         1651     :	result = 16'd255;
         1652     :	result = 16'd255;
         1653     :	result = 16'd255;
         1654     :	result = 16'd255;
         1655     :	result = 16'd255;
         1656     :	result = 16'd255;
         1657     :	result = 16'd255;
         1658     :	result = 16'd255;
         1659     :	result = 16'd255;
         1660     :	result = 16'd255;
         1661     :	result = 16'd255;
         1662     :	result = 16'd255;
         1663     :	result = 16'd255;
         1664     :	result = 16'd255;
         1665     :	result = 16'd255;
         1666     :	result = 16'd255;
         1667     :	result = 16'd255;
         1668     :	result = 16'd255;
         1669     :	result = 16'd255;
         1670     :	result = 16'd255;
         1671     :	result = 16'd255;
         1672     :	result = 16'd255;
         1673     :	result = 16'd255;
         1674     :	result = 16'd255;
         1675     :	result = 16'd255;
         1676     :	result = 16'd255;
         1677     :	result = 16'd255;
         1678     :	result = 16'd255;
         1679     :	result = 16'd255;
         1680     :	result = 16'd255;
         1681     :	result = 16'd255;
         1682     :	result = 16'd255;
         1683     :	result = 16'd255;
         1684     :	result = 16'd255;
         1685     :	result = 16'd255;
         1686     :	result = 16'd255;
         1687     :	result = 16'd255;
         1688     :	result = 16'd255;
         1689     :	result = 16'd255;
         1690     :	result = 16'd255;
         1691     :	result = 16'd255;
         1692     :	result = 16'd255;
         1693     :	result = 16'd255;
         1694     :	result = 16'd255;
         1695     :	result = 16'd255;
         1696     :	result = 16'd255;
         1697     :	result = 16'd255;
         1698     :	result = 16'd255;
         1699     :	result = 16'd255;
         1700     :	result = 16'd255;
         1701     :	result = 16'd255;
         1702     :	result = 16'd255;
         1703     :	result = 16'd255;
         1704     :	result = 16'd255;
         1705     :	result = 16'd255;
         1706     :	result = 16'd255;
         1707     :	result = 16'd255;
         1708     :	result = 16'd255;
         1709     :	result = 16'd255;
         1710     :	result = 16'd255;
         1711     :	result = 16'd255;
         1712     :	result = 16'd255;
         1713     :	result = 16'd255;
         1714     :	result = 16'd255;
         1715     :	result = 16'd255;
         1716     :	result = 16'd255;
         1717     :	result = 16'd255;
         1718     :	result = 16'd255;
         1719     :	result = 16'd255;
         1720     :	result = 16'd255;
         1721     :	result = 16'd255;
         1722     :	result = 16'd255;
         1723     :	result = 16'd255;
         1724     :	result = 16'd255;
         1725     :	result = 16'd255;
         1726     :	result = 16'd255;
         1727     :	result = 16'd255;
         1728     :	result = 16'd255;
         1729     :	result = 16'd255;
         1730     :	result = 16'd255;
         1731     :	result = 16'd255;
         1732     :	result = 16'd255;
         1733     :	result = 16'd255;
         1734     :	result = 16'd255;
         1735     :	result = 16'd255;
         1736     :	result = 16'd255;
         1737     :	result = 16'd255;
         1738     :	result = 16'd255;
         1739     :	result = 16'd255;
         1740     :	result = 16'd255;
         1741     :	result = 16'd255;
         1742     :	result = 16'd255;
         1743     :	result = 16'd255;
         1744     :	result = 16'd255;
         1745     :	result = 16'd255;
         1746     :	result = 16'd255;
         1747     :	result = 16'd255;
         1748     :	result = 16'd255;
         1749     :	result = 16'd255;
         1750     :	result = 16'd255;
         1751     :	result = 16'd255;
         1752     :	result = 16'd255;
         1753     :	result = 16'd255;
         1754     :	result = 16'd255;
         1755     :	result = 16'd255;
         1756     :	result = 16'd255;
         1757     :	result = 16'd255;
         1758     :	result = 16'd255;
         1759     :	result = 16'd255;
         1760     :	result = 16'd255;
         1761     :	result = 16'd255;
         1762     :	result = 16'd255;
         1763     :	result = 16'd255;
         1764     :	result = 16'd255;
         1765     :	result = 16'd255;
         1766     :	result = 16'd255;
         1767     :	result = 16'd255;
         1768     :	result = 16'd255;
         1769     :	result = 16'd255;
         1770     :	result = 16'd255;
         1771     :	result = 16'd255;
         1772     :	result = 16'd255;
         1773     :	result = 16'd255;
         1774     :	result = 16'd255;
         1775     :	result = 16'd255;
         1776     :	result = 16'd255;
         1777     :	result = 16'd255;
         1778     :	result = 16'd255;
         1779     :	result = 16'd255;
         1780     :	result = 16'd255;
         1781     :	result = 16'd255;
         1782     :	result = 16'd255;
         1783     :	result = 16'd255;
         1784     :	result = 16'd255;
         1785     :	result = 16'd255;
         1786     :	result = 16'd255;
         1787     :	result = 16'd255;
         1788     :	result = 16'd255;
         1789     :	result = 16'd255;
         1790     :	result = 16'd255;
         1791     :	result = 16'd255;

      endcase
   end

=======
//////////////////////////////////////////////////////////////////////////////////
// Engineer    : Achmad novel, Fauzan Ibrahim, Nicholas Teffandi
// Design Name : Autoencoder
// Module Name : sigmoid_lut
// Project Name: Autoencoder
//////////////////////////////////////////////////////////////////////////////////

// Input and Output is Unsigned

module sigmoid_lut {
   input wire [15:0] addr,
   output reg [15:0] addr
};

   always @(*) begin
      
      case (addr)
         63744    :	result = 16'd0
         63745    :	result = 16'd0
         63746    :	result = 16'd0
         63747    :	result = 16'd0
         63748    :	result = 16'd0
         63749    :	result = 16'd0
         63750    :	result = 16'd0
         63751    :	result = 16'd0
         63752    :	result = 16'd0
         63753    :	result = 16'd0
         63754    :	result = 16'd0
         63755    :	result = 16'd0
         63756    :	result = 16'd0
         63757    :	result = 16'd0
         63758    :	result = 16'd0
         63759    :	result = 16'd0
         63760    :	result = 16'd0
         63761    :	result = 16'd0
         63762    :	result = 16'd0
         63763    :	result = 16'd0
         63764    :	result = 16'd0
         63765    :	result = 16'd0
         63766    :	result = 16'd0
         63767    :	result = 16'd0
         63768    :	result = 16'd0
         63769    :	result = 16'd0
         63770    :	result = 16'd0
         63771    :	result = 16'd0
         63772    :	result = 16'd0
         63773    :	result = 16'd0
         63774    :	result = 16'd0
         63775    :	result = 16'd0
         63776    :	result = 16'd0
         63777    :	result = 16'd0
         63778    :	result = 16'd0
         63779    :	result = 16'd0
         63780    :	result = 16'd0
         63781    :	result = 16'd0
         63782    :	result = 16'd0
         63783    :	result = 16'd0
         63784    :	result = 16'd0
         63785    :	result = 16'd0
         63786    :	result = 16'd0
         63787    :	result = 16'd0
         63788    :	result = 16'd0
         63789    :	result = 16'd0
         63790    :	result = 16'd0
         63791    :	result = 16'd0
         63792    :	result = 16'd0
         63793    :	result = 16'd0
         63794    :	result = 16'd0
         63795    :	result = 16'd0
         63796    :	result = 16'd0
         63797    :	result = 16'd0
         63798    :	result = 16'd0
         63799    :	result = 16'd0
         63800    :	result = 16'd0
         63801    :	result = 16'd0
         63802    :	result = 16'd0
         63803    :	result = 16'd0
         63804    :	result = 16'd0
         63805    :	result = 16'd0
         63806    :	result = 16'd0
         63807    :	result = 16'd0
         63808    :	result = 16'd0
         63809    :	result = 16'd0
         63810    :	result = 16'd0
         63811    :	result = 16'd0
         63812    :	result = 16'd0
         63813    :	result = 16'd0
         63814    :	result = 16'd0
         63815    :	result = 16'd0
         63816    :	result = 16'd0
         63817    :	result = 16'd0
         63818    :	result = 16'd0
         63819    :	result = 16'd0
         63820    :	result = 16'd0
         63821    :	result = 16'd0
         63822    :	result = 16'd0
         63823    :	result = 16'd0
         63824    :	result = 16'd0
         63825    :	result = 16'd0
         63826    :	result = 16'd0
         63827    :	result = 16'd0
         63828    :	result = 16'd0
         63829    :	result = 16'd0
         63830    :	result = 16'd0
         63831    :	result = 16'd0
         63832    :	result = 16'd0
         63833    :	result = 16'd0
         63834    :	result = 16'd0
         63835    :	result = 16'd0
         63836    :	result = 16'd0
         63837    :	result = 16'd0
         63838    :	result = 16'd0
         63839    :	result = 16'd0
         63840    :	result = 16'd0
         63841    :	result = 16'd0
         63842    :	result = 16'd0
         63843    :	result = 16'd0
         63844    :	result = 16'd0
         63845    :	result = 16'd0
         63846    :	result = 16'd0
         63847    :	result = 16'd0
         63848    :	result = 16'd0
         63849    :	result = 16'd0
         63850    :	result = 16'd0
         63851    :	result = 16'd0
         63852    :	result = 16'd0
         63853    :	result = 16'd0
         63854    :	result = 16'd0
         63855    :	result = 16'd0
         63856    :	result = 16'd0
         63857    :	result = 16'd0
         63858    :	result = 16'd0
         63859    :	result = 16'd0
         63860    :	result = 16'd0
         63861    :	result = 16'd0
         63862    :	result = 16'd0
         63863    :	result = 16'd0
         63864    :	result = 16'd0
         63865    :	result = 16'd0
         63866    :	result = 16'd0
         63867    :	result = 16'd0
         63868    :	result = 16'd0
         63869    :	result = 16'd0
         63870    :	result = 16'd0
         63871    :	result = 16'd0
         63872    :	result = 16'd0
         63873    :	result = 16'd0
         63874    :	result = 16'd0
         63875    :	result = 16'd0
         63876    :	result = 16'd0
         63877    :	result = 16'd0
         63878    :	result = 16'd0
         63879    :	result = 16'd0
         63880    :	result = 16'd0
         63881    :	result = 16'd0
         63882    :	result = 16'd0
         63883    :	result = 16'd0
         63884    :	result = 16'd0
         63885    :	result = 16'd0
         63886    :	result = 16'd0
         63887    :	result = 16'd0
         63888    :	result = 16'd0
         63889    :	result = 16'd0
         63890    :	result = 16'd0
         63891    :	result = 16'd0
         63892    :	result = 16'd0
         63893    :	result = 16'd0
         63894    :	result = 16'd0
         63895    :	result = 16'd0
         63896    :	result = 16'd0
         63897    :	result = 16'd0
         63898    :	result = 16'd0
         63899    :	result = 16'd0
         63900    :	result = 16'd0
         63901    :	result = 16'd0
         63902    :	result = 16'd0
         63903    :	result = 16'd0
         63904    :	result = 16'd0
         63905    :	result = 16'd0
         63906    :	result = 16'd0
         63907    :	result = 16'd0
         63908    :	result = 16'd0
         63909    :	result = 16'd0
         63910    :	result = 16'd0
         63911    :	result = 16'd0
         63912    :	result = 16'd0
         63913    :	result = 16'd0
         63914    :	result = 16'd0
         63915    :	result = 16'd0
         63916    :	result = 16'd0
         63917    :	result = 16'd0
         63918    :	result = 16'd0
         63919    :	result = 16'd0
         63920    :	result = 16'd0
         63921    :	result = 16'd0
         63922    :	result = 16'd0
         63923    :	result = 16'd0
         63924    :	result = 16'd0
         63925    :	result = 16'd0
         63926    :	result = 16'd0
         63927    :	result = 16'd0
         63928    :	result = 16'd0
         63929    :	result = 16'd0
         63930    :	result = 16'd0
         63931    :	result = 16'd0
         63932    :	result = 16'd0
         63933    :	result = 16'd0
         63934    :	result = 16'd0
         63935    :	result = 16'd0
         63936    :	result = 16'd0
         63937    :	result = 16'd0
         63938    :	result = 16'd0
         63939    :	result = 16'd0
         63940    :	result = 16'd0
         63941    :	result = 16'd0
         63942    :	result = 16'd0
         63943    :	result = 16'd0
         63944    :	result = 16'd0
         63945    :	result = 16'd0
         63946    :	result = 16'd0
         63947    :	result = 16'd0
         63948    :	result = 16'd0
         63949    :	result = 16'd0
         63950    :	result = 16'd0
         63951    :	result = 16'd0
         63952    :	result = 16'd0
         63953    :	result = 16'd0
         63954    :	result = 16'd0
         63955    :	result = 16'd0
         63956    :	result = 16'd0
         63957    :	result = 16'd0
         63958    :	result = 16'd0
         63959    :	result = 16'd0
         63960    :	result = 16'd0
         63961    :	result = 16'd0
         63962    :	result = 16'd0
         63963    :	result = 16'd0
         63964    :	result = 16'd0
         63965    :	result = 16'd0
         63966    :	result = 16'd0
         63967    :	result = 16'd0
         63968    :	result = 16'd0
         63969    :	result = 16'd0
         63970    :	result = 16'd0
         63971    :	result = 16'd0
         63972    :	result = 16'd0
         63973    :	result = 16'd0
         63974    :	result = 16'd0
         63975    :	result = 16'd0
         63976    :	result = 16'd0
         63977    :	result = 16'd0
         63978    :	result = 16'd0
         63979    :	result = 16'd0
         63980    :	result = 16'd0
         63981    :	result = 16'd0
         63982    :	result = 16'd0
         63983    :	result = 16'd0
         63984    :	result = 16'd0
         63985    :	result = 16'd0
         63986    :	result = 16'd0
         63987    :	result = 16'd0
         63988    :	result = 16'd0
         63989    :	result = 16'd0
         63990    :	result = 16'd0
         63991    :	result = 16'd0
         63992    :	result = 16'd0
         63993    :	result = 16'd0
         63994    :	result = 16'd0
         63995    :	result = 16'd0
         63996    :	result = 16'd0
         63997    :	result = 16'd0
         63998    :	result = 16'd0
         63999    :	result = 16'd0
         64000    :	result = 16'd0
         64001    :	result = 16'd0
         64002    :	result = 16'd0
         64003    :	result = 16'd0
         64004    :	result = 16'd0
         64005    :	result = 16'd0
         64006    :	result = 16'd0
         64007    :	result = 16'd0
         64008    :	result = 16'd0
         64009    :	result = 16'd0
         64010    :	result = 16'd0
         64011    :	result = 16'd0
         64012    :	result = 16'd0
         64013    :	result = 16'd0
         64014    :	result = 16'd0
         64015    :	result = 16'd0
         64016    :	result = 16'd0
         64017    :	result = 16'd0
         64018    :	result = 16'd0
         64019    :	result = 16'd0
         64020    :	result = 16'd0
         64021    :	result = 16'd0
         64022    :	result = 16'd0
         64023    :	result = 16'd0
         64024    :	result = 16'd0
         64025    :	result = 16'd0
         64026    :	result = 16'd0
         64027    :	result = 16'd0
         64028    :	result = 16'd0
         64029    :	result = 16'd0
         64030    :	result = 16'd0
         64031    :	result = 16'd0
         64032    :	result = 16'd0
         64033    :	result = 16'd0
         64034    :	result = 16'd0
         64035    :	result = 16'd0
         64036    :	result = 16'd0
         64037    :	result = 16'd0
         64038    :	result = 16'd0
         64039    :	result = 16'd0
         64040    :	result = 16'd0
         64041    :	result = 16'd0
         64042    :	result = 16'd0
         64043    :	result = 16'd0
         64044    :	result = 16'd0
         64045    :	result = 16'd0
         64046    :	result = 16'd0
         64047    :	result = 16'd0
         64048    :	result = 16'd0
         64049    :	result = 16'd0
         64050    :	result = 16'd0
         64051    :	result = 16'd0
         64052    :	result = 16'd0
         64053    :	result = 16'd0
         64054    :	result = 16'd0
         64055    :	result = 16'd0
         64056    :	result = 16'd0
         64057    :	result = 16'd0
         64058    :	result = 16'd0
         64059    :	result = 16'd0
         64060    :	result = 16'd0
         64061    :	result = 16'd0
         64062    :	result = 16'd0
         64063    :	result = 16'd0
         64064    :	result = 16'd0
         64065    :	result = 16'd0
         64066    :	result = 16'd0
         64067    :	result = 16'd0
         64068    :	result = 16'd0
         64069    :	result = 16'd0
         64070    :	result = 16'd0
         64071    :	result = 16'd0
         64072    :	result = 16'd0
         64073    :	result = 16'd0
         64074    :	result = 16'd0
         64075    :	result = 16'd0
         64076    :	result = 16'd0
         64077    :	result = 16'd0
         64078    :	result = 16'd0
         64079    :	result = 16'd0
         64080    :	result = 16'd0
         64081    :	result = 16'd0
         64082    :	result = 16'd0
         64083    :	result = 16'd0
         64084    :	result = 16'd0
         64085    :	result = 16'd0
         64086    :	result = 16'd0
         64087    :	result = 16'd0
         64088    :	result = 16'd0
         64089    :	result = 16'd0
         64090    :	result = 16'd0
         64091    :	result = 16'd0
         64092    :	result = 16'd0
         64093    :	result = 16'd0
         64094    :	result = 16'd0
         64095    :	result = 16'd0
         64096    :	result = 16'd0
         64097    :	result = 16'd0
         64098    :	result = 16'd0
         64099    :	result = 16'd0
         64100    :	result = 16'd0
         64101    :	result = 16'd0
         64102    :	result = 16'd0
         64103    :	result = 16'd0
         64104    :	result = 16'd0
         64105    :	result = 16'd0
         64106    :	result = 16'd0
         64107    :	result = 16'd0
         64108    :	result = 16'd0
         64109    :	result = 16'd0
         64110    :	result = 16'd0
         64111    :	result = 16'd0
         64112    :	result = 16'd0
         64113    :	result = 16'd0
         64114    :	result = 16'd0
         64115    :	result = 16'd0
         64116    :	result = 16'd0
         64117    :	result = 16'd1
         64118    :	result = 16'd1
         64119    :	result = 16'd1
         64120    :	result = 16'd1
         64121    :	result = 16'd1
         64122    :	result = 16'd1
         64123    :	result = 16'd1
         64124    :	result = 16'd1
         64125    :	result = 16'd1
         64126    :	result = 16'd1
         64127    :	result = 16'd1
         64128    :	result = 16'd1
         64129    :	result = 16'd1
         64130    :	result = 16'd1
         64131    :	result = 16'd1
         64132    :	result = 16'd1
         64133    :	result = 16'd1
         64134    :	result = 16'd1
         64135    :	result = 16'd1
         64136    :	result = 16'd1
         64137    :	result = 16'd1
         64138    :	result = 16'd1
         64139    :	result = 16'd1
         64140    :	result = 16'd1
         64141    :	result = 16'd1
         64142    :	result = 16'd1
         64143    :	result = 16'd1
         64144    :	result = 16'd1
         64145    :	result = 16'd1
         64146    :	result = 16'd1
         64147    :	result = 16'd1
         64148    :	result = 16'd1
         64149    :	result = 16'd1
         64150    :	result = 16'd1
         64151    :	result = 16'd1
         64152    :	result = 16'd1
         64153    :	result = 16'd1
         64154    :	result = 16'd1
         64155    :	result = 16'd1
         64156    :	result = 16'd1
         64157    :	result = 16'd1
         64158    :	result = 16'd1
         64159    :	result = 16'd1
         64160    :	result = 16'd1
         64161    :	result = 16'd1
         64162    :	result = 16'd1
         64163    :	result = 16'd1
         64164    :	result = 16'd1
         64165    :	result = 16'd1
         64166    :	result = 16'd1
         64167    :	result = 16'd1
         64168    :	result = 16'd1
         64169    :	result = 16'd1
         64170    :	result = 16'd1
         64171    :	result = 16'd1
         64172    :	result = 16'd1
         64173    :	result = 16'd1
         64174    :	result = 16'd1
         64175    :	result = 16'd1
         64176    :	result = 16'd1
         64177    :	result = 16'd1
         64178    :	result = 16'd1
         64179    :	result = 16'd1
         64180    :	result = 16'd1
         64181    :	result = 16'd1
         64182    :	result = 16'd1
         64183    :	result = 16'd1
         64184    :	result = 16'd1
         64185    :	result = 16'd1
         64186    :	result = 16'd1
         64187    :	result = 16'd1
         64188    :	result = 16'd1
         64189    :	result = 16'd1
         64190    :	result = 16'd1
         64191    :	result = 16'd1
         64192    :	result = 16'd1
         64193    :	result = 16'd1
         64194    :	result = 16'd1
         64195    :	result = 16'd1
         64196    :	result = 16'd1
         64197    :	result = 16'd1
         64198    :	result = 16'd1
         64199    :	result = 16'd1
         64200    :	result = 16'd1
         64201    :	result = 16'd1
         64202    :	result = 16'd1
         64203    :	result = 16'd1
         64204    :	result = 16'd1
         64205    :	result = 16'd1
         64206    :	result = 16'd1
         64207    :	result = 16'd1
         64208    :	result = 16'd1
         64209    :	result = 16'd1
         64210    :	result = 16'd1
         64211    :	result = 16'd1
         64212    :	result = 16'd1
         64213    :	result = 16'd1
         64214    :	result = 16'd1
         64215    :	result = 16'd1
         64216    :	result = 16'd1
         64217    :	result = 16'd1
         64218    :	result = 16'd1
         64219    :	result = 16'd1
         64220    :	result = 16'd1
         64221    :	result = 16'd1
         64222    :	result = 16'd1
         64223    :	result = 16'd1
         64224    :	result = 16'd1
         64225    :	result = 16'd1
         64226    :	result = 16'd1
         64227    :	result = 16'd1
         64228    :	result = 16'd1
         64229    :	result = 16'd1
         64230    :	result = 16'd1
         64231    :	result = 16'd1
         64232    :	result = 16'd1
         64233    :	result = 16'd1
         64234    :	result = 16'd1
         64235    :	result = 16'd1
         64236    :	result = 16'd1
         64237    :	result = 16'd1
         64238    :	result = 16'd1
         64239    :	result = 16'd1
         64240    :	result = 16'd1
         64241    :	result = 16'd1
         64242    :	result = 16'd1
         64243    :	result = 16'd1
         64244    :	result = 16'd1
         64245    :	result = 16'd1
         64246    :	result = 16'd1
         64247    :	result = 16'd1
         64248    :	result = 16'd1
         64249    :	result = 16'd1
         64250    :	result = 16'd1
         64251    :	result = 16'd1
         64252    :	result = 16'd1
         64253    :	result = 16'd1
         64254    :	result = 16'd1
         64255    :	result = 16'd1
         64256    :	result = 16'd1
         64257    :	result = 16'd1
         64258    :	result = 16'd1
         64259    :	result = 16'd1
         64260    :	result = 16'd1
         64261    :	result = 16'd1
         64262    :	result = 16'd1
         64263    :	result = 16'd1
         64264    :	result = 16'd1
         64265    :	result = 16'd1
         64266    :	result = 16'd1
         64267    :	result = 16'd1
         64268    :	result = 16'd1
         64269    :	result = 16'd1
         64270    :	result = 16'd1
         64271    :	result = 16'd1
         64272    :	result = 16'd1
         64273    :	result = 16'd1
         64274    :	result = 16'd1
         64275    :	result = 16'd1
         64276    :	result = 16'd1
         64277    :	result = 16'd1
         64278    :	result = 16'd1
         64279    :	result = 16'd1
         64280    :	result = 16'd1
         64281    :	result = 16'd1
         64282    :	result = 16'd1
         64283    :	result = 16'd1
         64284    :	result = 16'd1
         64285    :	result = 16'd1
         64286    :	result = 16'd1
         64287    :	result = 16'd1
         64288    :	result = 16'd1
         64289    :	result = 16'd1
         64290    :	result = 16'd1
         64291    :	result = 16'd1
         64292    :	result = 16'd1
         64293    :	result = 16'd1
         64294    :	result = 16'd1
         64295    :	result = 16'd2
         64296    :	result = 16'd2
         64297    :	result = 16'd2
         64298    :	result = 16'd2
         64299    :	result = 16'd2
         64300    :	result = 16'd2
         64301    :	result = 16'd2
         64302    :	result = 16'd2
         64303    :	result = 16'd2
         64304    :	result = 16'd2
         64305    :	result = 16'd2
         64306    :	result = 16'd2
         64307    :	result = 16'd2
         64308    :	result = 16'd2
         64309    :	result = 16'd2
         64310    :	result = 16'd2
         64311    :	result = 16'd2
         64312    :	result = 16'd2
         64313    :	result = 16'd2
         64314    :	result = 16'd2
         64315    :	result = 16'd2
         64316    :	result = 16'd2
         64317    :	result = 16'd2
         64318    :	result = 16'd2
         64319    :	result = 16'd2
         64320    :	result = 16'd2
         64321    :	result = 16'd2
         64322    :	result = 16'd2
         64323    :	result = 16'd2
         64324    :	result = 16'd2
         64325    :	result = 16'd2
         64326    :	result = 16'd2
         64327    :	result = 16'd2
         64328    :	result = 16'd2
         64329    :	result = 16'd2
         64330    :	result = 16'd2
         64331    :	result = 16'd2
         64332    :	result = 16'd2
         64333    :	result = 16'd2
         64334    :	result = 16'd2
         64335    :	result = 16'd2
         64336    :	result = 16'd2
         64337    :	result = 16'd2
         64338    :	result = 16'd2
         64339    :	result = 16'd2
         64340    :	result = 16'd2
         64341    :	result = 16'd2
         64342    :	result = 16'd2
         64343    :	result = 16'd2
         64344    :	result = 16'd2
         64345    :	result = 16'd2
         64346    :	result = 16'd2
         64347    :	result = 16'd2
         64348    :	result = 16'd2
         64349    :	result = 16'd2
         64350    :	result = 16'd2
         64351    :	result = 16'd2
         64352    :	result = 16'd2
         64353    :	result = 16'd2
         64354    :	result = 16'd2
         64355    :	result = 16'd2
         64356    :	result = 16'd2
         64357    :	result = 16'd2
         64358    :	result = 16'd2
         64359    :	result = 16'd2
         64360    :	result = 16'd2
         64361    :	result = 16'd2
         64362    :	result = 16'd2
         64363    :	result = 16'd2
         64364    :	result = 16'd2
         64365    :	result = 16'd2
         64366    :	result = 16'd2
         64367    :	result = 16'd2
         64368    :	result = 16'd2
         64369    :	result = 16'd2
         64370    :	result = 16'd2
         64371    :	result = 16'd2
         64372    :	result = 16'd2
         64373    :	result = 16'd2
         64374    :	result = 16'd2
         64375    :	result = 16'd2
         64376    :	result = 16'd2
         64377    :	result = 16'd2
         64378    :	result = 16'd2
         64379    :	result = 16'd2
         64380    :	result = 16'd2
         64381    :	result = 16'd2
         64382    :	result = 16'd2
         64383    :	result = 16'd2
         64384    :	result = 16'd2
         64385    :	result = 16'd2
         64386    :	result = 16'd2
         64387    :	result = 16'd2
         64388    :	result = 16'd2
         64389    :	result = 16'd2
         64390    :	result = 16'd2
         64391    :	result = 16'd2
         64392    :	result = 16'd2
         64393    :	result = 16'd2
         64394    :	result = 16'd2
         64395    :	result = 16'd2
         64396    :	result = 16'd2
         64397    :	result = 16'd2
         64398    :	result = 16'd2
         64399    :	result = 16'd2
         64400    :	result = 16'd3
         64401    :	result = 16'd3
         64402    :	result = 16'd3
         64403    :	result = 16'd3
         64404    :	result = 16'd3
         64405    :	result = 16'd3
         64406    :	result = 16'd3
         64407    :	result = 16'd3
         64408    :	result = 16'd3
         64409    :	result = 16'd3
         64410    :	result = 16'd3
         64411    :	result = 16'd3
         64412    :	result = 16'd3
         64413    :	result = 16'd3
         64414    :	result = 16'd3
         64415    :	result = 16'd3
         64416    :	result = 16'd3
         64417    :	result = 16'd3
         64418    :	result = 16'd3
         64419    :	result = 16'd3
         64420    :	result = 16'd3
         64421    :	result = 16'd3
         64422    :	result = 16'd3
         64423    :	result = 16'd3
         64424    :	result = 16'd3
         64425    :	result = 16'd3
         64426    :	result = 16'd3
         64427    :	result = 16'd3
         64428    :	result = 16'd3
         64429    :	result = 16'd3
         64430    :	result = 16'd3
         64431    :	result = 16'd3
         64432    :	result = 16'd3
         64433    :	result = 16'd3
         64434    :	result = 16'd3
         64435    :	result = 16'd3
         64436    :	result = 16'd3
         64437    :	result = 16'd3
         64438    :	result = 16'd3
         64439    :	result = 16'd3
         64440    :	result = 16'd3
         64441    :	result = 16'd3
         64442    :	result = 16'd3
         64443    :	result = 16'd3
         64444    :	result = 16'd3
         64445    :	result = 16'd3
         64446    :	result = 16'd3
         64447    :	result = 16'd3
         64448    :	result = 16'd3
         64449    :	result = 16'd3
         64450    :	result = 16'd3
         64451    :	result = 16'd3
         64452    :	result = 16'd3
         64453    :	result = 16'd3
         64454    :	result = 16'd3
         64455    :	result = 16'd3
         64456    :	result = 16'd3
         64457    :	result = 16'd3
         64458    :	result = 16'd3
         64459    :	result = 16'd3
         64460    :	result = 16'd3
         64461    :	result = 16'd3
         64462    :	result = 16'd3
         64463    :	result = 16'd3
         64464    :	result = 16'd3
         64465    :	result = 16'd3
         64466    :	result = 16'd3
         64467    :	result = 16'd3
         64468    :	result = 16'd3
         64469    :	result = 16'd3
         64470    :	result = 16'd3
         64471    :	result = 16'd3
         64472    :	result = 16'd3
         64473    :	result = 16'd3
         64474    :	result = 16'd3
         64475    :	result = 16'd4
         64476    :	result = 16'd4
         64477    :	result = 16'd4
         64478    :	result = 16'd4
         64479    :	result = 16'd4
         64480    :	result = 16'd4
         64481    :	result = 16'd4
         64482    :	result = 16'd4
         64483    :	result = 16'd4
         64484    :	result = 16'd4
         64485    :	result = 16'd4
         64486    :	result = 16'd4
         64487    :	result = 16'd4
         64488    :	result = 16'd4
         64489    :	result = 16'd4
         64490    :	result = 16'd4
         64491    :	result = 16'd4
         64492    :	result = 16'd4
         64493    :	result = 16'd4
         64494    :	result = 16'd4
         64495    :	result = 16'd4
         64496    :	result = 16'd4
         64497    :	result = 16'd4
         64498    :	result = 16'd4
         64499    :	result = 16'd4
         64500    :	result = 16'd4
         64501    :	result = 16'd4
         64502    :	result = 16'd4
         64503    :	result = 16'd4
         64504    :	result = 16'd4
         64505    :	result = 16'd4
         64506    :	result = 16'd4
         64507    :	result = 16'd4
         64508    :	result = 16'd4
         64509    :	result = 16'd4
         64510    :	result = 16'd4
         64511    :	result = 16'd4
         64512    :	result = 16'd4
         64513    :	result = 16'd4
         64514    :	result = 16'd4
         64515    :	result = 16'd4
         64516    :	result = 16'd4
         64517    :	result = 16'd4
         64518    :	result = 16'd4
         64519    :	result = 16'd4
         64520    :	result = 16'd4
         64521    :	result = 16'd4
         64522    :	result = 16'd4
         64523    :	result = 16'd4
         64524    :	result = 16'd4
         64525    :	result = 16'd4
         64526    :	result = 16'd4
         64527    :	result = 16'd4
         64528    :	result = 16'd4
         64529    :	result = 16'd4
         64530    :	result = 16'd4
         64531    :	result = 16'd4
         64532    :	result = 16'd4
         64533    :	result = 16'd5
         64534    :	result = 16'd5
         64535    :	result = 16'd5
         64536    :	result = 16'd5
         64537    :	result = 16'd5
         64538    :	result = 16'd5
         64539    :	result = 16'd5
         64540    :	result = 16'd5
         64541    :	result = 16'd5
         64542    :	result = 16'd5
         64543    :	result = 16'd5
         64544    :	result = 16'd5
         64545    :	result = 16'd5
         64546    :	result = 16'd5
         64547    :	result = 16'd5
         64548    :	result = 16'd5
         64549    :	result = 16'd5
         64550    :	result = 16'd5
         64551    :	result = 16'd5
         64552    :	result = 16'd5
         64553    :	result = 16'd5
         64554    :	result = 16'd5
         64555    :	result = 16'd5
         64556    :	result = 16'd5
         64557    :	result = 16'd5
         64558    :	result = 16'd5
         64559    :	result = 16'd5
         64560    :	result = 16'd5
         64561    :	result = 16'd5
         64562    :	result = 16'd5
         64563    :	result = 16'd5
         64564    :	result = 16'd5
         64565    :	result = 16'd5
         64566    :	result = 16'd5
         64567    :	result = 16'd5
         64568    :	result = 16'd5
         64569    :	result = 16'd5
         64570    :	result = 16'd5
         64571    :	result = 16'd5
         64572    :	result = 16'd5
         64573    :	result = 16'd5
         64574    :	result = 16'd5
         64575    :	result = 16'd5
         64576    :	result = 16'd5
         64577    :	result = 16'd5
         64578    :	result = 16'd5
         64579    :	result = 16'd5
         64580    :	result = 16'd5
         64581    :	result = 16'd6
         64582    :	result = 16'd6
         64583    :	result = 16'd6
         64584    :	result = 16'd6
         64585    :	result = 16'd6
         64586    :	result = 16'd6
         64587    :	result = 16'd6
         64588    :	result = 16'd6
         64589    :	result = 16'd6
         64590    :	result = 16'd6
         64591    :	result = 16'd6
         64592    :	result = 16'd6
         64593    :	result = 16'd6
         64594    :	result = 16'd6
         64595    :	result = 16'd6
         64596    :	result = 16'd6
         64597    :	result = 16'd6
         64598    :	result = 16'd6
         64599    :	result = 16'd6
         64600    :	result = 16'd6
         64601    :	result = 16'd6
         64602    :	result = 16'd6
         64603    :	result = 16'd6
         64604    :	result = 16'd6
         64605    :	result = 16'd6
         64606    :	result = 16'd6
         64607    :	result = 16'd6
         64608    :	result = 16'd6
         64609    :	result = 16'd6
         64610    :	result = 16'd6
         64611    :	result = 16'd6
         64612    :	result = 16'd6
         64613    :	result = 16'd6
         64614    :	result = 16'd6
         64615    :	result = 16'd6
         64616    :	result = 16'd6
         64617    :	result = 16'd6
         64618    :	result = 16'd6
         64619    :	result = 16'd6
         64620    :	result = 16'd6
         64621    :	result = 16'd7
         64622    :	result = 16'd7
         64623    :	result = 16'd7
         64624    :	result = 16'd7
         64625    :	result = 16'd7
         64626    :	result = 16'd7
         64627    :	result = 16'd7
         64628    :	result = 16'd7
         64629    :	result = 16'd7
         64630    :	result = 16'd7
         64631    :	result = 16'd7
         64632    :	result = 16'd7
         64633    :	result = 16'd7
         64634    :	result = 16'd7
         64635    :	result = 16'd7
         64636    :	result = 16'd7
         64637    :	result = 16'd7
         64638    :	result = 16'd7
         64639    :	result = 16'd7
         64640    :	result = 16'd7
         64641    :	result = 16'd7
         64642    :	result = 16'd7
         64643    :	result = 16'd7
         64644    :	result = 16'd7
         64645    :	result = 16'd7
         64646    :	result = 16'd7
         64647    :	result = 16'd7
         64648    :	result = 16'd7
         64649    :	result = 16'd7
         64650    :	result = 16'd7
         64651    :	result = 16'd7
         64652    :	result = 16'd7
         64653    :	result = 16'd7
         64654    :	result = 16'd7
         64655    :	result = 16'd7
         64656    :	result = 16'd8
         64657    :	result = 16'd8
         64658    :	result = 16'd8
         64659    :	result = 16'd8
         64660    :	result = 16'd8
         64661    :	result = 16'd8
         64662    :	result = 16'd8
         64663    :	result = 16'd8
         64664    :	result = 16'd8
         64665    :	result = 16'd8
         64666    :	result = 16'd8
         64667    :	result = 16'd8
         64668    :	result = 16'd8
         64669    :	result = 16'd8
         64670    :	result = 16'd8
         64671    :	result = 16'd8
         64672    :	result = 16'd8
         64673    :	result = 16'd8
         64674    :	result = 16'd8
         64675    :	result = 16'd8
         64676    :	result = 16'd8
         64677    :	result = 16'd8
         64678    :	result = 16'd8
         64679    :	result = 16'd8
         64680    :	result = 16'd8
         64681    :	result = 16'd8
         64682    :	result = 16'd8
         64683    :	result = 16'd8
         64684    :	result = 16'd8
         64685    :	result = 16'd8
         64686    :	result = 16'd8
         64687    :	result = 16'd8
         64688    :	result = 16'd9
         64689    :	result = 16'd9
         64690    :	result = 16'd9
         64691    :	result = 16'd9
         64692    :	result = 16'd9
         64693    :	result = 16'd9
         64694    :	result = 16'd9
         64695    :	result = 16'd9
         64696    :	result = 16'd9
         64697    :	result = 16'd9
         64698    :	result = 16'd9
         64699    :	result = 16'd9
         64700    :	result = 16'd9
         64701    :	result = 16'd9
         64702    :	result = 16'd9
         64703    :	result = 16'd9
         64704    :	result = 16'd9
         64705    :	result = 16'd9
         64706    :	result = 16'd9
         64707    :	result = 16'd9
         64708    :	result = 16'd9
         64709    :	result = 16'd9
         64710    :	result = 16'd9
         64711    :	result = 16'd9
         64712    :	result = 16'd9
         64713    :	result = 16'd9
         64714    :	result = 16'd9
         64715    :	result = 16'd9
         64716    :	result = 16'd10
         64717    :	result = 16'd10
         64718    :	result = 16'd10
         64719    :	result = 16'd10
         64720    :	result = 16'd10
         64721    :	result = 16'd10
         64722    :	result = 16'd10
         64723    :	result = 16'd10
         64724    :	result = 16'd10
         64725    :	result = 16'd10
         64726    :	result = 16'd10
         64727    :	result = 16'd10
         64728    :	result = 16'd10
         64729    :	result = 16'd10
         64730    :	result = 16'd10
         64731    :	result = 16'd10
         64732    :	result = 16'd10
         64733    :	result = 16'd10
         64734    :	result = 16'd10
         64735    :	result = 16'd10
         64736    :	result = 16'd10
         64737    :	result = 16'd10
         64738    :	result = 16'd10
         64739    :	result = 16'd10
         64740    :	result = 16'd10
         64741    :	result = 16'd11
         64742    :	result = 16'd11
         64743    :	result = 16'd11
         64744    :	result = 16'd11
         64745    :	result = 16'd11
         64746    :	result = 16'd11
         64747    :	result = 16'd11
         64748    :	result = 16'd11
         64749    :	result = 16'd11
         64750    :	result = 16'd11
         64751    :	result = 16'd11
         64752    :	result = 16'd11
         64753    :	result = 16'd11
         64754    :	result = 16'd11
         64755    :	result = 16'd11
         64756    :	result = 16'd11
         64757    :	result = 16'd11
         64758    :	result = 16'd11
         64759    :	result = 16'd11
         64760    :	result = 16'd11
         64761    :	result = 16'd11
         64762    :	result = 16'd11
         64763    :	result = 16'd11
         64764    :	result = 16'd12
         64765    :	result = 16'd12
         64766    :	result = 16'd12
         64767    :	result = 16'd12
         64768    :	result = 16'd12
         64769    :	result = 16'd12
         64770    :	result = 16'd12
         64771    :	result = 16'd12
         64772    :	result = 16'd12
         64773    :	result = 16'd12
         64774    :	result = 16'd12
         64775    :	result = 16'd12
         64776    :	result = 16'd12
         64777    :	result = 16'd12
         64778    :	result = 16'd12
         64779    :	result = 16'd12
         64780    :	result = 16'd12
         64781    :	result = 16'd12
         64782    :	result = 16'd12
         64783    :	result = 16'd12
         64784    :	result = 16'd12
         64785    :	result = 16'd12
         64786    :	result = 16'd13
         64787    :	result = 16'd13
         64788    :	result = 16'd13
         64789    :	result = 16'd13
         64790    :	result = 16'd13
         64791    :	result = 16'd13
         64792    :	result = 16'd13
         64793    :	result = 16'd13
         64794    :	result = 16'd13
         64795    :	result = 16'd13
         64796    :	result = 16'd13
         64797    :	result = 16'd13
         64798    :	result = 16'd13
         64799    :	result = 16'd13
         64800    :	result = 16'd13
         64801    :	result = 16'd13
         64802    :	result = 16'd13
         64803    :	result = 16'd13
         64804    :	result = 16'd13
         64805    :	result = 16'd13
         64806    :	result = 16'd14
         64807    :	result = 16'd14
         64808    :	result = 16'd14
         64809    :	result = 16'd14
         64810    :	result = 16'd14
         64811    :	result = 16'd14
         64812    :	result = 16'd14
         64813    :	result = 16'd14
         64814    :	result = 16'd14
         64815    :	result = 16'd14
         64816    :	result = 16'd14
         64817    :	result = 16'd14
         64818    :	result = 16'd14
         64819    :	result = 16'd14
         64820    :	result = 16'd14
         64821    :	result = 16'd14
         64822    :	result = 16'd14
         64823    :	result = 16'd14
         64824    :	result = 16'd14
         64825    :	result = 16'd15
         64826    :	result = 16'd15
         64827    :	result = 16'd15
         64828    :	result = 16'd15
         64829    :	result = 16'd15
         64830    :	result = 16'd15
         64831    :	result = 16'd15
         64832    :	result = 16'd15
         64833    :	result = 16'd15
         64834    :	result = 16'd15
         64835    :	result = 16'd15
         64836    :	result = 16'd15
         64837    :	result = 16'd15
         64838    :	result = 16'd15
         64839    :	result = 16'd15
         64840    :	result = 16'd15
         64841    :	result = 16'd15
         64842    :	result = 16'd16
         64843    :	result = 16'd16
         64844    :	result = 16'd16
         64845    :	result = 16'd16
         64846    :	result = 16'd16
         64847    :	result = 16'd16
         64848    :	result = 16'd16
         64849    :	result = 16'd16
         64850    :	result = 16'd16
         64851    :	result = 16'd16
         64852    :	result = 16'd16
         64853    :	result = 16'd16
         64854    :	result = 16'd16
         64855    :	result = 16'd16
         64856    :	result = 16'd16
         64857    :	result = 16'd16
         64858    :	result = 16'd16
         64859    :	result = 16'd17
         64860    :	result = 16'd17
         64861    :	result = 16'd17
         64862    :	result = 16'd17
         64863    :	result = 16'd17
         64864    :	result = 16'd17
         64865    :	result = 16'd17
         64866    :	result = 16'd17
         64867    :	result = 16'd17
         64868    :	result = 16'd17
         64869    :	result = 16'd17
         64870    :	result = 16'd17
         64871    :	result = 16'd17
         64872    :	result = 16'd17
         64873    :	result = 16'd17
         64874    :	result = 16'd17
         64875    :	result = 16'd18
         64876    :	result = 16'd18
         64877    :	result = 16'd18
         64878    :	result = 16'd18
         64879    :	result = 16'd18
         64880    :	result = 16'd18
         64881    :	result = 16'd18
         64882    :	result = 16'd18
         64883    :	result = 16'd18
         64884    :	result = 16'd18
         64885    :	result = 16'd18
         64886    :	result = 16'd18
         64887    :	result = 16'd18
         64888    :	result = 16'd18
         64889    :	result = 16'd19
         64890    :	result = 16'd19
         64891    :	result = 16'd19
         64892    :	result = 16'd19
         64893    :	result = 16'd19
         64894    :	result = 16'd19
         64895    :	result = 16'd19
         64896    :	result = 16'd19
         64897    :	result = 16'd19
         64898    :	result = 16'd19
         64899    :	result = 16'd19
         64900    :	result = 16'd19
         64901    :	result = 16'd19
         64902    :	result = 16'd19
         64903    :	result = 16'd19
         64904    :	result = 16'd20
         64905    :	result = 16'd20
         64906    :	result = 16'd20
         64907    :	result = 16'd20
         64908    :	result = 16'd20
         64909    :	result = 16'd20
         64910    :	result = 16'd20
         64911    :	result = 16'd20
         64912    :	result = 16'd20
         64913    :	result = 16'd20
         64914    :	result = 16'd20
         64915    :	result = 16'd20
         64916    :	result = 16'd20
         64917    :	result = 16'd21
         64918    :	result = 16'd21
         64919    :	result = 16'd21
         64920    :	result = 16'd21
         64921    :	result = 16'd21
         64922    :	result = 16'd21
         64923    :	result = 16'd21
         64924    :	result = 16'd21
         64925    :	result = 16'd21
         64926    :	result = 16'd21
         64927    :	result = 16'd21
         64928    :	result = 16'd21
         64929    :	result = 16'd21
         64930    :	result = 16'd22
         64931    :	result = 16'd22
         64932    :	result = 16'd22
         64933    :	result = 16'd22
         64934    :	result = 16'd22
         64935    :	result = 16'd22
         64936    :	result = 16'd22
         64937    :	result = 16'd22
         64938    :	result = 16'd22
         64939    :	result = 16'd22
         64940    :	result = 16'd22
         64941    :	result = 16'd22
         64942    :	result = 16'd22
         64943    :	result = 16'd23
         64944    :	result = 16'd23
         64945    :	result = 16'd23
         64946    :	result = 16'd23
         64947    :	result = 16'd23
         64948    :	result = 16'd23
         64949    :	result = 16'd23
         64950    :	result = 16'd23
         64951    :	result = 16'd23
         64952    :	result = 16'd23
         64953    :	result = 16'd23
         64954    :	result = 16'd23
         64955    :	result = 16'd24
         64956    :	result = 16'd24
         64957    :	result = 16'd24
         64958    :	result = 16'd24
         64959    :	result = 16'd24
         64960    :	result = 16'd24
         64961    :	result = 16'd24
         64962    :	result = 16'd24
         64963    :	result = 16'd24
         64964    :	result = 16'd24
         64965    :	result = 16'd24
         64966    :	result = 16'd25
         64967    :	result = 16'd25
         64968    :	result = 16'd25
         64969    :	result = 16'd25
         64970    :	result = 16'd25
         64971    :	result = 16'd25
         64972    :	result = 16'd25
         64973    :	result = 16'd25
         64974    :	result = 16'd25
         64975    :	result = 16'd25
         64976    :	result = 16'd25
         64977    :	result = 16'd26
         64978    :	result = 16'd26
         64979    :	result = 16'd26
         64980    :	result = 16'd26
         64981    :	result = 16'd26
         64982    :	result = 16'd26
         64983    :	result = 16'd26
         64984    :	result = 16'd26
         64985    :	result = 16'd26
         64986    :	result = 16'd26
         64987    :	result = 16'd26
         64988    :	result = 16'd27
         64989    :	result = 16'd27
         64990    :	result = 16'd27
         64991    :	result = 16'd27
         64992    :	result = 16'd27
         64993    :	result = 16'd27
         64994    :	result = 16'd27
         64995    :	result = 16'd27
         64996    :	result = 16'd27
         64997    :	result = 16'd27
         64998    :	result = 16'd27
         64999    :	result = 16'd28
         65000    :	result = 16'd28
         65001    :	result = 16'd28
         65002    :	result = 16'd28
         65003    :	result = 16'd28
         65004    :	result = 16'd28
         65005    :	result = 16'd28
         65006    :	result = 16'd28
         65007    :	result = 16'd28
         65008    :	result = 16'd28
         65009    :	result = 16'd29
         65010    :	result = 16'd29
         65011    :	result = 16'd29
         65012    :	result = 16'd29
         65013    :	result = 16'd29
         65014    :	result = 16'd29
         65015    :	result = 16'd29
         65016    :	result = 16'd29
         65017    :	result = 16'd29
         65018    :	result = 16'd29
         65019    :	result = 16'd30
         65020    :	result = 16'd30
         65021    :	result = 16'd30
         65022    :	result = 16'd30
         65023    :	result = 16'd30
         65024    :	result = 16'd30
         65025    :	result = 16'd30
         65026    :	result = 16'd30
         65027    :	result = 16'd30
         65028    :	result = 16'd31
         65029    :	result = 16'd31
         65030    :	result = 16'd31
         65031    :	result = 16'd31
         65032    :	result = 16'd31
         65033    :	result = 16'd31
         65034    :	result = 16'd31
         65035    :	result = 16'd31
         65036    :	result = 16'd31
         65037    :	result = 16'd32
         65038    :	result = 16'd32
         65039    :	result = 16'd32
         65040    :	result = 16'd32
         65041    :	result = 16'd32
         65042    :	result = 16'd32
         65043    :	result = 16'd32
         65044    :	result = 16'd32
         65045    :	result = 16'd32
         65046    :	result = 16'd33
         65047    :	result = 16'd33
         65048    :	result = 16'd33
         65049    :	result = 16'd33
         65050    :	result = 16'd33
         65051    :	result = 16'd33
         65052    :	result = 16'd33
         65053    :	result = 16'd33
         65054    :	result = 16'd33
         65055    :	result = 16'd34
         65056    :	result = 16'd34
         65057    :	result = 16'd34
         65058    :	result = 16'd34
         65059    :	result = 16'd34
         65060    :	result = 16'd34
         65061    :	result = 16'd34
         65062    :	result = 16'd34
         65063    :	result = 16'd34
         65064    :	result = 16'd35
         65065    :	result = 16'd35
         65066    :	result = 16'd35
         65067    :	result = 16'd35
         65068    :	result = 16'd35
         65069    :	result = 16'd35
         65070    :	result = 16'd35
         65071    :	result = 16'd35
         65072    :	result = 16'd36
         65073    :	result = 16'd36
         65074    :	result = 16'd36
         65075    :	result = 16'd36
         65076    :	result = 16'd36
         65077    :	result = 16'd36
         65078    :	result = 16'd36
         65079    :	result = 16'd36
         65080    :	result = 16'd37
         65081    :	result = 16'd37
         65082    :	result = 16'd37
         65083    :	result = 16'd37
         65084    :	result = 16'd37
         65085    :	result = 16'd37
         65086    :	result = 16'd37
         65087    :	result = 16'd37
         65088    :	result = 16'd38
         65089    :	result = 16'd38
         65090    :	result = 16'd38
         65091    :	result = 16'd38
         65092    :	result = 16'd38
         65093    :	result = 16'd38
         65094    :	result = 16'd38
         65095    :	result = 16'd38
         65096    :	result = 16'd39
         65097    :	result = 16'd39
         65098    :	result = 16'd39
         65099    :	result = 16'd39
         65100    :	result = 16'd39
         65101    :	result = 16'd39
         65102    :	result = 16'd39
         65103    :	result = 16'd39
         65104    :	result = 16'd40
         65105    :	result = 16'd40
         65106    :	result = 16'd40
         65107    :	result = 16'd40
         65108    :	result = 16'd40
         65109    :	result = 16'd40
         65110    :	result = 16'd40
         65111    :	result = 16'd41
         65112    :	result = 16'd41
         65113    :	result = 16'd41
         65114    :	result = 16'd41
         65115    :	result = 16'd41
         65116    :	result = 16'd41
         65117    :	result = 16'd41
         65118    :	result = 16'd41
         65119    :	result = 16'd42
         65120    :	result = 16'd42
         65121    :	result = 16'd42
         65122    :	result = 16'd42
         65123    :	result = 16'd42
         65124    :	result = 16'd42
         65125    :	result = 16'd42
         65126    :	result = 16'd43
         65127    :	result = 16'd43
         65128    :	result = 16'd43
         65129    :	result = 16'd43
         65130    :	result = 16'd43
         65131    :	result = 16'd43
         65132    :	result = 16'd43
         65133    :	result = 16'd44
         65134    :	result = 16'd44
         65135    :	result = 16'd44
         65136    :	result = 16'd44
         65137    :	result = 16'd44
         65138    :	result = 16'd44
         65139    :	result = 16'd44
         65140    :	result = 16'd45
         65141    :	result = 16'd45
         65142    :	result = 16'd45
         65143    :	result = 16'd45
         65144    :	result = 16'd45
         65145    :	result = 16'd45
         65146    :	result = 16'd45
         65147    :	result = 16'd46
         65148    :	result = 16'd46
         65149    :	result = 16'd46
         65150    :	result = 16'd46
         65151    :	result = 16'd46
         65152    :	result = 16'd46
         65153    :	result = 16'd46
         65154    :	result = 16'd47
         65155    :	result = 16'd47
         65156    :	result = 16'd47
         65157    :	result = 16'd47
         65158    :	result = 16'd47
         65159    :	result = 16'd47
         65160    :	result = 16'd48
         65161    :	result = 16'd48
         65162    :	result = 16'd48
         65163    :	result = 16'd48
         65164    :	result = 16'd48
         65165    :	result = 16'd48
         65166    :	result = 16'd48
         65167    :	result = 16'd49
         65168    :	result = 16'd49
         65169    :	result = 16'd49
         65170    :	result = 16'd49
         65171    :	result = 16'd49
         65172    :	result = 16'd49
         65173    :	result = 16'd50
         65174    :	result = 16'd50
         65175    :	result = 16'd50
         65176    :	result = 16'd50
         65177    :	result = 16'd50
         65178    :	result = 16'd50
         65179    :	result = 16'd51
         65180    :	result = 16'd51
         65181    :	result = 16'd51
         65182    :	result = 16'd51
         65183    :	result = 16'd51
         65184    :	result = 16'd51
         65185    :	result = 16'd51
         65186    :	result = 16'd52
         65187    :	result = 16'd52
         65188    :	result = 16'd52
         65189    :	result = 16'd52
         65190    :	result = 16'd52
         65191    :	result = 16'd52
         65192    :	result = 16'd53
         65193    :	result = 16'd53
         65194    :	result = 16'd53
         65195    :	result = 16'd53
         65196    :	result = 16'd53
         65197    :	result = 16'd53
         65198    :	result = 16'd54
         65199    :	result = 16'd54
         65200    :	result = 16'd54
         65201    :	result = 16'd54
         65202    :	result = 16'd54
         65203    :	result = 16'd54
         65204    :	result = 16'd55
         65205    :	result = 16'd55
         65206    :	result = 16'd55
         65207    :	result = 16'd55
         65208    :	result = 16'd55
         65209    :	result = 16'd55
         65210    :	result = 16'd56
         65211    :	result = 16'd56
         65212    :	result = 16'd56
         65213    :	result = 16'd56
         65214    :	result = 16'd56
         65215    :	result = 16'd57
         65216    :	result = 16'd57
         65217    :	result = 16'd57
         65218    :	result = 16'd57
         65219    :	result = 16'd57
         65220    :	result = 16'd57
         65221    :	result = 16'd58
         65222    :	result = 16'd58
         65223    :	result = 16'd58
         65224    :	result = 16'd58
         65225    :	result = 16'd58
         65226    :	result = 16'd58
         65227    :	result = 16'd59
         65228    :	result = 16'd59
         65229    :	result = 16'd59
         65230    :	result = 16'd59
         65231    :	result = 16'd59
         65232    :	result = 16'd60
         65233    :	result = 16'd60
         65234    :	result = 16'd60
         65235    :	result = 16'd60
         65236    :	result = 16'd60
         65237    :	result = 16'd60
         65238    :	result = 16'd61
         65239    :	result = 16'd61
         65240    :	result = 16'd61
         65241    :	result = 16'd61
         65242    :	result = 16'd61
         65243    :	result = 16'd62
         65244    :	result = 16'd62
         65245    :	result = 16'd62
         65246    :	result = 16'd62
         65247    :	result = 16'd62
         65248    :	result = 16'd62
         65249    :	result = 16'd63
         65250    :	result = 16'd63
         65251    :	result = 16'd63
         65252    :	result = 16'd63
         65253    :	result = 16'd63
         65254    :	result = 16'd64
         65255    :	result = 16'd64
         65256    :	result = 16'd64
         65257    :	result = 16'd64
         65258    :	result = 16'd64
         65259    :	result = 16'd64
         65260    :	result = 16'd65
         65261    :	result = 16'd65
         65262    :	result = 16'd65
         65263    :	result = 16'd65
         65264    :	result = 16'd65
         65265    :	result = 16'd66
         65266    :	result = 16'd66
         65267    :	result = 16'd66
         65268    :	result = 16'd66
         65269    :	result = 16'd66
         65270    :	result = 16'd67
         65271    :	result = 16'd67
         65272    :	result = 16'd67
         65273    :	result = 16'd67
         65274    :	result = 16'd67
         65275    :	result = 16'd68
         65276    :	result = 16'd68
         65277    :	result = 16'd68
         65278    :	result = 16'd68
         65279    :	result = 16'd68
         65280    :	result = 16'd69
         65281    :	result = 16'd69
         65282    :	result = 16'd69
         65283    :	result = 16'd69
         65284    :	result = 16'd69
         65285    :	result = 16'd70
         65286    :	result = 16'd70
         65287    :	result = 16'd70
         65288    :	result = 16'd70
         65289    :	result = 16'd70
         65290    :	result = 16'd71
         65291    :	result = 16'd71
         65292    :	result = 16'd71
         65293    :	result = 16'd71
         65294    :	result = 16'd71
         65295    :	result = 16'd72
         65296    :	result = 16'd72
         65297    :	result = 16'd72
         65298    :	result = 16'd72
         65299    :	result = 16'd72
         65300    :	result = 16'd73
         65301    :	result = 16'd73
         65302    :	result = 16'd73
         65303    :	result = 16'd73
         65304    :	result = 16'd73
         65305    :	result = 16'd74
         65306    :	result = 16'd74
         65307    :	result = 16'd74
         65308    :	result = 16'd74
         65309    :	result = 16'd74
         65310    :	result = 16'd75
         65311    :	result = 16'd75
         65312    :	result = 16'd75
         65313    :	result = 16'd75
         65314    :	result = 16'd75
         65315    :	result = 16'd76
         65316    :	result = 16'd76
         65317    :	result = 16'd76
         65318    :	result = 16'd76
         65319    :	result = 16'd76
         65320    :	result = 16'd77
         65321    :	result = 16'd77
         65322    :	result = 16'd77
         65323    :	result = 16'd77
         65324    :	result = 16'd78
         65325    :	result = 16'd78
         65326    :	result = 16'd78
         65327    :	result = 16'd78
         65328    :	result = 16'd78
         65329    :	result = 16'd79
         65330    :	result = 16'd79
         65331    :	result = 16'd79
         65332    :	result = 16'd79
         65333    :	result = 16'd79
         65334    :	result = 16'd80
         65335    :	result = 16'd80
         65336    :	result = 16'd80
         65337    :	result = 16'd80
         65338    :	result = 16'd81
         65339    :	result = 16'd81
         65340    :	result = 16'd81
         65341    :	result = 16'd81
         65342    :	result = 16'd81
         65343    :	result = 16'd82
         65344    :	result = 16'd82
         65345    :	result = 16'd82
         65346    :	result = 16'd82
         65347    :	result = 16'd83
         65348    :	result = 16'd83
         65349    :	result = 16'd83
         65350    :	result = 16'd83
         65351    :	result = 16'd83
         65352    :	result = 16'd84
         65353    :	result = 16'd84
         65354    :	result = 16'd84
         65355    :	result = 16'd84
         65356    :	result = 16'd84
         65357    :	result = 16'd85
         65358    :	result = 16'd85
         65359    :	result = 16'd85
         65360    :	result = 16'd85
         65361    :	result = 16'd86
         65362    :	result = 16'd86
         65363    :	result = 16'd86
         65364    :	result = 16'd86
         65365    :	result = 16'd86
         65366    :	result = 16'd87
         65367    :	result = 16'd87
         65368    :	result = 16'd87
         65369    :	result = 16'd87
         65370    :	result = 16'd88
         65371    :	result = 16'd88
         65372    :	result = 16'd88
         65373    :	result = 16'd88
         65374    :	result = 16'd89
         65375    :	result = 16'd89
         65376    :	result = 16'd89
         65377    :	result = 16'd89
         65378    :	result = 16'd89
         65379    :	result = 16'd90
         65380    :	result = 16'd90
         65381    :	result = 16'd90
         65382    :	result = 16'd90
         65383    :	result = 16'd91
         65384    :	result = 16'd91
         65385    :	result = 16'd91
         65386    :	result = 16'd91
         65387    :	result = 16'd91
         65388    :	result = 16'd92
         65389    :	result = 16'd92
         65390    :	result = 16'd92
         65391    :	result = 16'd92
         65392    :	result = 16'd93
         65393    :	result = 16'd93
         65394    :	result = 16'd93
         65395    :	result = 16'd93
         65396    :	result = 16'd94
         65397    :	result = 16'd94
         65398    :	result = 16'd94
         65399    :	result = 16'd94
         65400    :	result = 16'd95
         65401    :	result = 16'd95
         65402    :	result = 16'd95
         65403    :	result = 16'd95
         65404    :	result = 16'd95
         65405    :	result = 16'd96
         65406    :	result = 16'd96
         65407    :	result = 16'd96
         65408    :	result = 16'd96
         65409    :	result = 16'd97
         65410    :	result = 16'd97
         65411    :	result = 16'd97
         65412    :	result = 16'd97
         65413    :	result = 16'd98
         65414    :	result = 16'd98
         65415    :	result = 16'd98
         65416    :	result = 16'd98
         65417    :	result = 16'd99
         65418    :	result = 16'd99
         65419    :	result = 16'd99
         65420    :	result = 16'd99
         65421    :	result = 16'd99
         65422    :	result = 16'd100
         65423    :	result = 16'd100
         65424    :	result = 16'd100
         65425    :	result = 16'd100
         65426    :	result = 16'd101
         65427    :	result = 16'd101
         65428    :	result = 16'd101
         65429    :	result = 16'd101
         65430    :	result = 16'd102
         65431    :	result = 16'd102
         65432    :	result = 16'd102
         65433    :	result = 16'd102
         65434    :	result = 16'd103
         65435    :	result = 16'd103
         65436    :	result = 16'd103
         65437    :	result = 16'd103
         65438    :	result = 16'd104
         65439    :	result = 16'd104
         65440    :	result = 16'd104
         65441    :	result = 16'd104
         65442    :	result = 16'd105
         65443    :	result = 16'd105
         65444    :	result = 16'd105
         65445    :	result = 16'd105
         65446    :	result = 16'd105
         65447    :	result = 16'd106
         65448    :	result = 16'd106
         65449    :	result = 16'd106
         65450    :	result = 16'd106
         65451    :	result = 16'd107
         65452    :	result = 16'd107
         65453    :	result = 16'd107
         65454    :	result = 16'd107
         65455    :	result = 16'd108
         65456    :	result = 16'd108
         65457    :	result = 16'd108
         65458    :	result = 16'd108
         65459    :	result = 16'd109
         65460    :	result = 16'd109
         65461    :	result = 16'd109
         65462    :	result = 16'd109
         65463    :	result = 16'd110
         65464    :	result = 16'd110
         65465    :	result = 16'd110
         65466    :	result = 16'd110
         65467    :	result = 16'd111
         65468    :	result = 16'd111
         65469    :	result = 16'd111
         65470    :	result = 16'd111
         65471    :	result = 16'd112
         65472    :	result = 16'd112
         65473    :	result = 16'd112
         65474    :	result = 16'd112
         65475    :	result = 16'd113
         65476    :	result = 16'd113
         65477    :	result = 16'd113
         65478    :	result = 16'd113
         65479    :	result = 16'd114
         65480    :	result = 16'd114
         65481    :	result = 16'd114
         65482    :	result = 16'd114
         65483    :	result = 16'd115
         65484    :	result = 16'd115
         65485    :	result = 16'd115
         65486    :	result = 16'd115
         65487    :	result = 16'd116
         65488    :	result = 16'd116
         65489    :	result = 16'd116
         65490    :	result = 16'd116
         65491    :	result = 16'd117
         65492    :	result = 16'd117
         65493    :	result = 16'd117
         65494    :	result = 16'd117
         65495    :	result = 16'd118
         65496    :	result = 16'd118
         65497    :	result = 16'd118
         65498    :	result = 16'd118
         65499    :	result = 16'd119
         65500    :	result = 16'd119
         65501    :	result = 16'd119
         65502    :	result = 16'd119
         65503    :	result = 16'd120
         65504    :	result = 16'd120
         65505    :	result = 16'd120
         65506    :	result = 16'd120
         65507    :	result = 16'd121
         65508    :	result = 16'd121
         65509    :	result = 16'd121
         65510    :	result = 16'd121
         65511    :	result = 16'd122
         65512    :	result = 16'd122
         65513    :	result = 16'd122
         65514    :	result = 16'd122
         65515    :	result = 16'd123
         65516    :	result = 16'd123
         65517    :	result = 16'd123
         65518    :	result = 16'd123
         65519    :	result = 16'd124
         65520    :	result = 16'd124
         65521    :	result = 16'd124
         65522    :	result = 16'd124
         65523    :	result = 16'd125
         65524    :	result = 16'd125
         65525    :	result = 16'd125
         65526    :	result = 16'd125
         65527    :	result = 16'd126
         65528    :	result = 16'd126
         65529    :	result = 16'd126
         65530    :	result = 16'd126
         65531    :	result = 16'd127
         65532    :	result = 16'd127
         65533    :	result = 16'd127
         65534    :	result = 16'd127
         65535    :	result = 16'd128
         0        :	result = 16'd128
         1        :	result = 16'd128
         2        :	result = 16'd128
         3        :	result = 16'd128
         4        :	result = 16'd129
         5        :	result = 16'd129
         6        :	result = 16'd129
         7        :	result = 16'd129
         8        :	result = 16'd130
         9        :	result = 16'd130
         10       :	result = 16'd130
         11       :	result = 16'd130
         12       :	result = 16'd131
         13       :	result = 16'd131
         14       :	result = 16'd131
         15       :	result = 16'd131
         16       :	result = 16'd132
         17       :	result = 16'd132
         18       :	result = 16'd132
         19       :	result = 16'd132
         20       :	result = 16'd133
         21       :	result = 16'd133
         22       :	result = 16'd133
         23       :	result = 16'd133
         24       :	result = 16'd134
         25       :	result = 16'd134
         26       :	result = 16'd134
         27       :	result = 16'd134
         28       :	result = 16'd135
         29       :	result = 16'd135
         30       :	result = 16'd135
         31       :	result = 16'd135
         32       :	result = 16'd136
         33       :	result = 16'd136
         34       :	result = 16'd136
         35       :	result = 16'd136
         36       :	result = 16'd137
         37       :	result = 16'd137
         38       :	result = 16'd137
         39       :	result = 16'd137
         40       :	result = 16'd138
         41       :	result = 16'd138
         42       :	result = 16'd138
         43       :	result = 16'd138
         44       :	result = 16'd139
         45       :	result = 16'd139
         46       :	result = 16'd139
         47       :	result = 16'd139
         48       :	result = 16'd140
         49       :	result = 16'd140
         50       :	result = 16'd140
         51       :	result = 16'd140
         52       :	result = 16'd141
         53       :	result = 16'd141
         54       :	result = 16'd141
         55       :	result = 16'd141
         56       :	result = 16'd142
         57       :	result = 16'd142
         58       :	result = 16'd142
         59       :	result = 16'd142
         60       :	result = 16'd143
         61       :	result = 16'd143
         62       :	result = 16'd143
         63       :	result = 16'd143
         64       :	result = 16'd144
         65       :	result = 16'd144
         66       :	result = 16'd144
         67       :	result = 16'd144
         68       :	result = 16'd145
         69       :	result = 16'd145
         70       :	result = 16'd145
         71       :	result = 16'd145
         72       :	result = 16'd146
         73       :	result = 16'd146
         74       :	result = 16'd146
         75       :	result = 16'd146
         76       :	result = 16'd147
         77       :	result = 16'd147
         78       :	result = 16'd147
         79       :	result = 16'd147
         80       :	result = 16'd148
         81       :	result = 16'd148
         82       :	result = 16'd148
         83       :	result = 16'd148
         84       :	result = 16'd149
         85       :	result = 16'd149
         86       :	result = 16'd149
         87       :	result = 16'd149
         88       :	result = 16'd150
         89       :	result = 16'd150
         90       :	result = 16'd150
         91       :	result = 16'd150
         92       :	result = 16'd150
         93       :	result = 16'd151
         94       :	result = 16'd151
         95       :	result = 16'd151
         96       :	result = 16'd151
         97       :	result = 16'd152
         98       :	result = 16'd152
         99       :	result = 16'd152
         100      :	result = 16'd152
         101      :	result = 16'd153
         102      :	result = 16'd153
         103      :	result = 16'd153
         104      :	result = 16'd153
         105      :	result = 16'd154
         106      :	result = 16'd154
         107      :	result = 16'd154
         108      :	result = 16'd154
         109      :	result = 16'd155
         110      :	result = 16'd155
         111      :	result = 16'd155
         112      :	result = 16'd155
         113      :	result = 16'd156
         114      :	result = 16'd156
         115      :	result = 16'd156
         116      :	result = 16'd156
         117      :	result = 16'd156
         118      :	result = 16'd157
         119      :	result = 16'd157
         120      :	result = 16'd157
         121      :	result = 16'd157
         122      :	result = 16'd158
         123      :	result = 16'd158
         124      :	result = 16'd158
         125      :	result = 16'd158
         126      :	result = 16'd159
         127      :	result = 16'd159
         128      :	result = 16'd159
         129      :	result = 16'd159
         130      :	result = 16'd160
         131      :	result = 16'd160
         132      :	result = 16'd160
         133      :	result = 16'd160
         134      :	result = 16'd160
         135      :	result = 16'd161
         136      :	result = 16'd161
         137      :	result = 16'd161
         138      :	result = 16'd161
         139      :	result = 16'd162
         140      :	result = 16'd162
         141      :	result = 16'd162
         142      :	result = 16'd162
         143      :	result = 16'd163
         144      :	result = 16'd163
         145      :	result = 16'd163
         146      :	result = 16'd163
         147      :	result = 16'd164
         148      :	result = 16'd164
         149      :	result = 16'd164
         150      :	result = 16'd164
         151      :	result = 16'd164
         152      :	result = 16'd165
         153      :	result = 16'd165
         154      :	result = 16'd165
         155      :	result = 16'd165
         156      :	result = 16'd166
         157      :	result = 16'd166
         158      :	result = 16'd166
         159      :	result = 16'd166
         160      :	result = 16'd166
         161      :	result = 16'd167
         162      :	result = 16'd167
         163      :	result = 16'd167
         164      :	result = 16'd167
         165      :	result = 16'd168
         166      :	result = 16'd168
         167      :	result = 16'd168
         168      :	result = 16'd168
         169      :	result = 16'd169
         170      :	result = 16'd169
         171      :	result = 16'd169
         172      :	result = 16'd169
         173      :	result = 16'd169
         174      :	result = 16'd170
         175      :	result = 16'd170
         176      :	result = 16'd170
         177      :	result = 16'd170
         178      :	result = 16'd171
         179      :	result = 16'd171
         180      :	result = 16'd171
         181      :	result = 16'd171
         182      :	result = 16'd171
         183      :	result = 16'd172
         184      :	result = 16'd172
         185      :	result = 16'd172
         186      :	result = 16'd172
         187      :	result = 16'd172
         188      :	result = 16'd173
         189      :	result = 16'd173
         190      :	result = 16'd173
         191      :	result = 16'd173
         192      :	result = 16'd174
         193      :	result = 16'd174
         194      :	result = 16'd174
         195      :	result = 16'd174
         196      :	result = 16'd174
         197      :	result = 16'd175
         198      :	result = 16'd175
         199      :	result = 16'd175
         200      :	result = 16'd175
         201      :	result = 16'd176
         202      :	result = 16'd176
         203      :	result = 16'd176
         204      :	result = 16'd176
         205      :	result = 16'd176
         206      :	result = 16'd177
         207      :	result = 16'd177
         208      :	result = 16'd177
         209      :	result = 16'd177
         210      :	result = 16'd177
         211      :	result = 16'd178
         212      :	result = 16'd178
         213      :	result = 16'd178
         214      :	result = 16'd178
         215      :	result = 16'd179
         216      :	result = 16'd179
         217      :	result = 16'd179
         218      :	result = 16'd179
         219      :	result = 16'd179
         220      :	result = 16'd180
         221      :	result = 16'd180
         222      :	result = 16'd180
         223      :	result = 16'd180
         224      :	result = 16'd180
         225      :	result = 16'd181
         226      :	result = 16'd181
         227      :	result = 16'd181
         228      :	result = 16'd181
         229      :	result = 16'd181
         230      :	result = 16'd182
         231      :	result = 16'd182
         232      :	result = 16'd182
         233      :	result = 16'd182
         234      :	result = 16'd182
         235      :	result = 16'd183
         236      :	result = 16'd183
         237      :	result = 16'd183
         238      :	result = 16'd183
         239      :	result = 16'd183
         240      :	result = 16'd184
         241      :	result = 16'd184
         242      :	result = 16'd184
         243      :	result = 16'd184
         244      :	result = 16'd184
         245      :	result = 16'd185
         246      :	result = 16'd185
         247      :	result = 16'd185
         248      :	result = 16'd185
         249      :	result = 16'd185
         250      :	result = 16'd186
         251      :	result = 16'd186
         252      :	result = 16'd186
         253      :	result = 16'd186
         254      :	result = 16'd186
         255      :	result = 16'd187
         256      :	result = 16'd187
         257      :	result = 16'd187
         258      :	result = 16'd187
         259      :	result = 16'd187
         260      :	result = 16'd188
         261      :	result = 16'd188
         262      :	result = 16'd188
         263      :	result = 16'd188
         264      :	result = 16'd188
         265      :	result = 16'd189
         266      :	result = 16'd189
         267      :	result = 16'd189
         268      :	result = 16'd189
         269      :	result = 16'd189
         270      :	result = 16'd190
         271      :	result = 16'd190
         272      :	result = 16'd190
         273      :	result = 16'd190
         274      :	result = 16'd190
         275      :	result = 16'd191
         276      :	result = 16'd191
         277      :	result = 16'd191
         278      :	result = 16'd191
         279      :	result = 16'd191
         280      :	result = 16'd191
         281      :	result = 16'd192
         282      :	result = 16'd192
         283      :	result = 16'd192
         284      :	result = 16'd192
         285      :	result = 16'd192
         286      :	result = 16'd193
         287      :	result = 16'd193
         288      :	result = 16'd193
         289      :	result = 16'd193
         290      :	result = 16'd193
         291      :	result = 16'd193
         292      :	result = 16'd194
         293      :	result = 16'd194
         294      :	result = 16'd194
         295      :	result = 16'd194
         296      :	result = 16'd194
         297      :	result = 16'd195
         298      :	result = 16'd195
         299      :	result = 16'd195
         300      :	result = 16'd195
         301      :	result = 16'd195
         302      :	result = 16'd195
         303      :	result = 16'd196
         304      :	result = 16'd196
         305      :	result = 16'd196
         306      :	result = 16'd196
         307      :	result = 16'd196
         308      :	result = 16'd197
         309      :	result = 16'd197
         310      :	result = 16'd197
         311      :	result = 16'd197
         312      :	result = 16'd197
         313      :	result = 16'd197
         314      :	result = 16'd198
         315      :	result = 16'd198
         316      :	result = 16'd198
         317      :	result = 16'd198
         318      :	result = 16'd198
         319      :	result = 16'd198
         320      :	result = 16'd199
         321      :	result = 16'd199
         322      :	result = 16'd199
         323      :	result = 16'd199
         324      :	result = 16'd199
         325      :	result = 16'd200
         326      :	result = 16'd200
         327      :	result = 16'd200
         328      :	result = 16'd200
         329      :	result = 16'd200
         330      :	result = 16'd200
         331      :	result = 16'd201
         332      :	result = 16'd201
         333      :	result = 16'd201
         334      :	result = 16'd201
         335      :	result = 16'd201
         336      :	result = 16'd201
         337      :	result = 16'd202
         338      :	result = 16'd202
         339      :	result = 16'd202
         340      :	result = 16'd202
         341      :	result = 16'd202
         342      :	result = 16'd202
         343      :	result = 16'd203
         344      :	result = 16'd203
         345      :	result = 16'd203
         346      :	result = 16'd203
         347      :	result = 16'd203
         348      :	result = 16'd203
         349      :	result = 16'd204
         350      :	result = 16'd204
         351      :	result = 16'd204
         352      :	result = 16'd204
         353      :	result = 16'd204
         354      :	result = 16'd204
         355      :	result = 16'd204
         356      :	result = 16'd205
         357      :	result = 16'd205
         358      :	result = 16'd205
         359      :	result = 16'd205
         360      :	result = 16'd205
         361      :	result = 16'd205
         362      :	result = 16'd206
         363      :	result = 16'd206
         364      :	result = 16'd206
         365      :	result = 16'd206
         366      :	result = 16'd206
         367      :	result = 16'd206
         368      :	result = 16'd207
         369      :	result = 16'd207
         370      :	result = 16'd207
         371      :	result = 16'd207
         372      :	result = 16'd207
         373      :	result = 16'd207
         374      :	result = 16'd207
         375      :	result = 16'd208
         376      :	result = 16'd208
         377      :	result = 16'd208
         378      :	result = 16'd208
         379      :	result = 16'd208
         380      :	result = 16'd208
         381      :	result = 16'd209
         382      :	result = 16'd209
         383      :	result = 16'd209
         384      :	result = 16'd209
         385      :	result = 16'd209
         386      :	result = 16'd209
         387      :	result = 16'd209
         388      :	result = 16'd210
         389      :	result = 16'd210
         390      :	result = 16'd210
         391      :	result = 16'd210
         392      :	result = 16'd210
         393      :	result = 16'd210
         394      :	result = 16'd210
         395      :	result = 16'd211
         396      :	result = 16'd211
         397      :	result = 16'd211
         398      :	result = 16'd211
         399      :	result = 16'd211
         400      :	result = 16'd211
         401      :	result = 16'd211
         402      :	result = 16'd212
         403      :	result = 16'd212
         404      :	result = 16'd212
         405      :	result = 16'd212
         406      :	result = 16'd212
         407      :	result = 16'd212
         408      :	result = 16'd212
         409      :	result = 16'd213
         410      :	result = 16'd213
         411      :	result = 16'd213
         412      :	result = 16'd213
         413      :	result = 16'd213
         414      :	result = 16'd213
         415      :	result = 16'd213
         416      :	result = 16'd214
         417      :	result = 16'd214
         418      :	result = 16'd214
         419      :	result = 16'd214
         420      :	result = 16'd214
         421      :	result = 16'd214
         422      :	result = 16'd214
         423      :	result = 16'd214
         424      :	result = 16'd215
         425      :	result = 16'd215
         426      :	result = 16'd215
         427      :	result = 16'd215
         428      :	result = 16'd215
         429      :	result = 16'd215
         430      :	result = 16'd215
         431      :	result = 16'd216
         432      :	result = 16'd216
         433      :	result = 16'd216
         434      :	result = 16'd216
         435      :	result = 16'd216
         436      :	result = 16'd216
         437      :	result = 16'd216
         438      :	result = 16'd216
         439      :	result = 16'd217
         440      :	result = 16'd217
         441      :	result = 16'd217
         442      :	result = 16'd217
         443      :	result = 16'd217
         444      :	result = 16'd217
         445      :	result = 16'd217
         446      :	result = 16'd217
         447      :	result = 16'd218
         448      :	result = 16'd218
         449      :	result = 16'd218
         450      :	result = 16'd218
         451      :	result = 16'd218
         452      :	result = 16'd218
         453      :	result = 16'd218
         454      :	result = 16'd218
         455      :	result = 16'd219
         456      :	result = 16'd219
         457      :	result = 16'd219
         458      :	result = 16'd219
         459      :	result = 16'd219
         460      :	result = 16'd219
         461      :	result = 16'd219
         462      :	result = 16'd219
         463      :	result = 16'd220
         464      :	result = 16'd220
         465      :	result = 16'd220
         466      :	result = 16'd220
         467      :	result = 16'd220
         468      :	result = 16'd220
         469      :	result = 16'd220
         470      :	result = 16'd220
         471      :	result = 16'd221
         472      :	result = 16'd221
         473      :	result = 16'd221
         474      :	result = 16'd221
         475      :	result = 16'd221
         476      :	result = 16'd221
         477      :	result = 16'd221
         478      :	result = 16'd221
         479      :	result = 16'd221
         480      :	result = 16'd222
         481      :	result = 16'd222
         482      :	result = 16'd222
         483      :	result = 16'd222
         484      :	result = 16'd222
         485      :	result = 16'd222
         486      :	result = 16'd222
         487      :	result = 16'd222
         488      :	result = 16'd222
         489      :	result = 16'd223
         490      :	result = 16'd223
         491      :	result = 16'd223
         492      :	result = 16'd223
         493      :	result = 16'd223
         494      :	result = 16'd223
         495      :	result = 16'd223
         496      :	result = 16'd223
         497      :	result = 16'd223
         498      :	result = 16'd224
         499      :	result = 16'd224
         500      :	result = 16'd224
         501      :	result = 16'd224
         502      :	result = 16'd224
         503      :	result = 16'd224
         504      :	result = 16'd224
         505      :	result = 16'd224
         506      :	result = 16'd224
         507      :	result = 16'd225
         508      :	result = 16'd225
         509      :	result = 16'd225
         510      :	result = 16'd225
         511      :	result = 16'd225
         512      :	result = 16'd225
         513      :	result = 16'd225
         514      :	result = 16'd225
         515      :	result = 16'd225
         516      :	result = 16'd226
         517      :	result = 16'd226
         518      :	result = 16'd226
         519      :	result = 16'd226
         520      :	result = 16'd226
         521      :	result = 16'd226
         522      :	result = 16'd226
         523      :	result = 16'd226
         524      :	result = 16'd226
         525      :	result = 16'd226
         526      :	result = 16'd227
         527      :	result = 16'd227
         528      :	result = 16'd227
         529      :	result = 16'd227
         530      :	result = 16'd227
         531      :	result = 16'd227
         532      :	result = 16'd227
         533      :	result = 16'd227
         534      :	result = 16'd227
         535      :	result = 16'd227
         536      :	result = 16'd228
         537      :	result = 16'd228
         538      :	result = 16'd228
         539      :	result = 16'd228
         540      :	result = 16'd228
         541      :	result = 16'd228
         542      :	result = 16'd228
         543      :	result = 16'd228
         544      :	result = 16'd228
         545      :	result = 16'd228
         546      :	result = 16'd228
         547      :	result = 16'd229
         548      :	result = 16'd229
         549      :	result = 16'd229
         550      :	result = 16'd229
         551      :	result = 16'd229
         552      :	result = 16'd229
         553      :	result = 16'd229
         554      :	result = 16'd229
         555      :	result = 16'd229
         556      :	result = 16'd229
         557      :	result = 16'd229
         558      :	result = 16'd230
         559      :	result = 16'd230
         560      :	result = 16'd230
         561      :	result = 16'd230
         562      :	result = 16'd230
         563      :	result = 16'd230
         564      :	result = 16'd230
         565      :	result = 16'd230
         566      :	result = 16'd230
         567      :	result = 16'd230
         568      :	result = 16'd230
         569      :	result = 16'd231
         570      :	result = 16'd231
         571      :	result = 16'd231
         572      :	result = 16'd231
         573      :	result = 16'd231
         574      :	result = 16'd231
         575      :	result = 16'd231
         576      :	result = 16'd231
         577      :	result = 16'd231
         578      :	result = 16'd231
         579      :	result = 16'd231
         580      :	result = 16'd232
         581      :	result = 16'd232
         582      :	result = 16'd232
         583      :	result = 16'd232
         584      :	result = 16'd232
         585      :	result = 16'd232
         586      :	result = 16'd232
         587      :	result = 16'd232
         588      :	result = 16'd232
         589      :	result = 16'd232
         590      :	result = 16'd232
         591      :	result = 16'd232
         592      :	result = 16'd233
         593      :	result = 16'd233
         594      :	result = 16'd233
         595      :	result = 16'd233
         596      :	result = 16'd233
         597      :	result = 16'd233
         598      :	result = 16'd233
         599      :	result = 16'd233
         600      :	result = 16'd233
         601      :	result = 16'd233
         602      :	result = 16'd233
         603      :	result = 16'd233
         604      :	result = 16'd233
         605      :	result = 16'd234
         606      :	result = 16'd234
         607      :	result = 16'd234
         608      :	result = 16'd234
         609      :	result = 16'd234
         610      :	result = 16'd234
         611      :	result = 16'd234
         612      :	result = 16'd234
         613      :	result = 16'd234
         614      :	result = 16'd234
         615      :	result = 16'd234
         616      :	result = 16'd234
         617      :	result = 16'd234
         618      :	result = 16'd235
         619      :	result = 16'd235
         620      :	result = 16'd235
         621      :	result = 16'd235
         622      :	result = 16'd235
         623      :	result = 16'd235
         624      :	result = 16'd235
         625      :	result = 16'd235
         626      :	result = 16'd235
         627      :	result = 16'd235
         628      :	result = 16'd235
         629      :	result = 16'd235
         630      :	result = 16'd235
         631      :	result = 16'd236
         632      :	result = 16'd236
         633      :	result = 16'd236
         634      :	result = 16'd236
         635      :	result = 16'd236
         636      :	result = 16'd236
         637      :	result = 16'd236
         638      :	result = 16'd236
         639      :	result = 16'd236
         640      :	result = 16'd236
         641      :	result = 16'd236
         642      :	result = 16'd236
         643      :	result = 16'd236
         644      :	result = 16'd236
         645      :	result = 16'd236
         646      :	result = 16'd237
         647      :	result = 16'd237
         648      :	result = 16'd237
         649      :	result = 16'd237
         650      :	result = 16'd237
         651      :	result = 16'd237
         652      :	result = 16'd237
         653      :	result = 16'd237
         654      :	result = 16'd237
         655      :	result = 16'd237
         656      :	result = 16'd237
         657      :	result = 16'd237
         658      :	result = 16'd237
         659      :	result = 16'd237
         660      :	result = 16'd238
         661      :	result = 16'd238
         662      :	result = 16'd238
         663      :	result = 16'd238
         664      :	result = 16'd238
         665      :	result = 16'd238
         666      :	result = 16'd238
         667      :	result = 16'd238
         668      :	result = 16'd238
         669      :	result = 16'd238
         670      :	result = 16'd238
         671      :	result = 16'd238
         672      :	result = 16'd238
         673      :	result = 16'd238
         674      :	result = 16'd238
         675      :	result = 16'd238
         676      :	result = 16'd239
         677      :	result = 16'd239
         678      :	result = 16'd239
         679      :	result = 16'd239
         680      :	result = 16'd239
         681      :	result = 16'd239
         682      :	result = 16'd239
         683      :	result = 16'd239
         684      :	result = 16'd239
         685      :	result = 16'd239
         686      :	result = 16'd239
         687      :	result = 16'd239
         688      :	result = 16'd239
         689      :	result = 16'd239
         690      :	result = 16'd239
         691      :	result = 16'd239
         692      :	result = 16'd239
         693      :	result = 16'd240
         694      :	result = 16'd240
         695      :	result = 16'd240
         696      :	result = 16'd240
         697      :	result = 16'd240
         698      :	result = 16'd240
         699      :	result = 16'd240
         700      :	result = 16'd240
         701      :	result = 16'd240
         702      :	result = 16'd240
         703      :	result = 16'd240
         704      :	result = 16'd240
         705      :	result = 16'd240
         706      :	result = 16'd240
         707      :	result = 16'd240
         708      :	result = 16'd240
         709      :	result = 16'd240
         710      :	result = 16'd241
         711      :	result = 16'd241
         712      :	result = 16'd241
         713      :	result = 16'd241
         714      :	result = 16'd241
         715      :	result = 16'd241
         716      :	result = 16'd241
         717      :	result = 16'd241
         718      :	result = 16'd241
         719      :	result = 16'd241
         720      :	result = 16'd241
         721      :	result = 16'd241
         722      :	result = 16'd241
         723      :	result = 16'd241
         724      :	result = 16'd241
         725      :	result = 16'd241
         726      :	result = 16'd241
         727      :	result = 16'd241
         728      :	result = 16'd241
         729      :	result = 16'd242
         730      :	result = 16'd242
         731      :	result = 16'd242
         732      :	result = 16'd242
         733      :	result = 16'd242
         734      :	result = 16'd242
         735      :	result = 16'd242
         736      :	result = 16'd242
         737      :	result = 16'd242
         738      :	result = 16'd242
         739      :	result = 16'd242
         740      :	result = 16'd242
         741      :	result = 16'd242
         742      :	result = 16'd242
         743      :	result = 16'd242
         744      :	result = 16'd242
         745      :	result = 16'd242
         746      :	result = 16'd242
         747      :	result = 16'd242
         748      :	result = 16'd242
         749      :	result = 16'd243
         750      :	result = 16'd243
         751      :	result = 16'd243
         752      :	result = 16'd243
         753      :	result = 16'd243
         754      :	result = 16'd243
         755      :	result = 16'd243
         756      :	result = 16'd243
         757      :	result = 16'd243
         758      :	result = 16'd243
         759      :	result = 16'd243
         760      :	result = 16'd243
         761      :	result = 16'd243
         762      :	result = 16'd243
         763      :	result = 16'd243
         764      :	result = 16'd243
         765      :	result = 16'd243
         766      :	result = 16'd243
         767      :	result = 16'd243
         768      :	result = 16'd243
         769      :	result = 16'd243
         770      :	result = 16'd243
         771      :	result = 16'd244
         772      :	result = 16'd244
         773      :	result = 16'd244
         774      :	result = 16'd244
         775      :	result = 16'd244
         776      :	result = 16'd244
         777      :	result = 16'd244
         778      :	result = 16'd244
         779      :	result = 16'd244
         780      :	result = 16'd244
         781      :	result = 16'd244
         782      :	result = 16'd244
         783      :	result = 16'd244
         784      :	result = 16'd244
         785      :	result = 16'd244
         786      :	result = 16'd244
         787      :	result = 16'd244
         788      :	result = 16'd244
         789      :	result = 16'd244
         790      :	result = 16'd244
         791      :	result = 16'd244
         792      :	result = 16'd244
         793      :	result = 16'd244
         794      :	result = 16'd245
         795      :	result = 16'd245
         796      :	result = 16'd245
         797      :	result = 16'd245
         798      :	result = 16'd245
         799      :	result = 16'd245
         800      :	result = 16'd245
         801      :	result = 16'd245
         802      :	result = 16'd245
         803      :	result = 16'd245
         804      :	result = 16'd245
         805      :	result = 16'd245
         806      :	result = 16'd245
         807      :	result = 16'd245
         808      :	result = 16'd245
         809      :	result = 16'd245
         810      :	result = 16'd245
         811      :	result = 16'd245
         812      :	result = 16'd245
         813      :	result = 16'd245
         814      :	result = 16'd245
         815      :	result = 16'd245
         816      :	result = 16'd245
         817      :	result = 16'd245
         818      :	result = 16'd245
         819      :	result = 16'd246
         820      :	result = 16'd246
         821      :	result = 16'd246
         822      :	result = 16'd246
         823      :	result = 16'd246
         824      :	result = 16'd246
         825      :	result = 16'd246
         826      :	result = 16'd246
         827      :	result = 16'd246
         828      :	result = 16'd246
         829      :	result = 16'd246
         830      :	result = 16'd246
         831      :	result = 16'd246
         832      :	result = 16'd246
         833      :	result = 16'd246
         834      :	result = 16'd246
         835      :	result = 16'd246
         836      :	result = 16'd246
         837      :	result = 16'd246
         838      :	result = 16'd246
         839      :	result = 16'd246
         840      :	result = 16'd246
         841      :	result = 16'd246
         842      :	result = 16'd246
         843      :	result = 16'd246
         844      :	result = 16'd246
         845      :	result = 16'd246
         846      :	result = 16'd246
         847      :	result = 16'd247
         848      :	result = 16'd247
         849      :	result = 16'd247
         850      :	result = 16'd247
         851      :	result = 16'd247
         852      :	result = 16'd247
         853      :	result = 16'd247
         854      :	result = 16'd247
         855      :	result = 16'd247
         856      :	result = 16'd247
         857      :	result = 16'd247
         858      :	result = 16'd247
         859      :	result = 16'd247
         860      :	result = 16'd247
         861      :	result = 16'd247
         862      :	result = 16'd247
         863      :	result = 16'd247
         864      :	result = 16'd247
         865      :	result = 16'd247
         866      :	result = 16'd247
         867      :	result = 16'd247
         868      :	result = 16'd247
         869      :	result = 16'd247
         870      :	result = 16'd247
         871      :	result = 16'd247
         872      :	result = 16'd247
         873      :	result = 16'd247
         874      :	result = 16'd247
         875      :	result = 16'd247
         876      :	result = 16'd247
         877      :	result = 16'd247
         878      :	result = 16'd247
         879      :	result = 16'd248
         880      :	result = 16'd248
         881      :	result = 16'd248
         882      :	result = 16'd248
         883      :	result = 16'd248
         884      :	result = 16'd248
         885      :	result = 16'd248
         886      :	result = 16'd248
         887      :	result = 16'd248
         888      :	result = 16'd248
         889      :	result = 16'd248
         890      :	result = 16'd248
         891      :	result = 16'd248
         892      :	result = 16'd248
         893      :	result = 16'd248
         894      :	result = 16'd248
         895      :	result = 16'd248
         896      :	result = 16'd248
         897      :	result = 16'd248
         898      :	result = 16'd248
         899      :	result = 16'd248
         900      :	result = 16'd248
         901      :	result = 16'd248
         902      :	result = 16'd248
         903      :	result = 16'd248
         904      :	result = 16'd248
         905      :	result = 16'd248
         906      :	result = 16'd248
         907      :	result = 16'd248
         908      :	result = 16'd248
         909      :	result = 16'd248
         910      :	result = 16'd248
         911      :	result = 16'd248
         912      :	result = 16'd248
         913      :	result = 16'd248
         914      :	result = 16'd249
         915      :	result = 16'd249
         916      :	result = 16'd249
         917      :	result = 16'd249
         918      :	result = 16'd249
         919      :	result = 16'd249
         920      :	result = 16'd249
         921      :	result = 16'd249
         922      :	result = 16'd249
         923      :	result = 16'd249
         924      :	result = 16'd249
         925      :	result = 16'd249
         926      :	result = 16'd249
         927      :	result = 16'd249
         928      :	result = 16'd249
         929      :	result = 16'd249
         930      :	result = 16'd249
         931      :	result = 16'd249
         932      :	result = 16'd249
         933      :	result = 16'd249
         934      :	result = 16'd249
         935      :	result = 16'd249
         936      :	result = 16'd249
         937      :	result = 16'd249
         938      :	result = 16'd249
         939      :	result = 16'd249
         940      :	result = 16'd249
         941      :	result = 16'd249
         942      :	result = 16'd249
         943      :	result = 16'd249
         944      :	result = 16'd249
         945      :	result = 16'd249
         946      :	result = 16'd249
         947      :	result = 16'd249
         948      :	result = 16'd249
         949      :	result = 16'd249
         950      :	result = 16'd249
         951      :	result = 16'd249
         952      :	result = 16'd249
         953      :	result = 16'd249
         954      :	result = 16'd250
         955      :	result = 16'd250
         956      :	result = 16'd250
         957      :	result = 16'd250
         958      :	result = 16'd250
         959      :	result = 16'd250
         960      :	result = 16'd250
         961      :	result = 16'd250
         962      :	result = 16'd250
         963      :	result = 16'd250
         964      :	result = 16'd250
         965      :	result = 16'd250
         966      :	result = 16'd250
         967      :	result = 16'd250
         968      :	result = 16'd250
         969      :	result = 16'd250
         970      :	result = 16'd250
         971      :	result = 16'd250
         972      :	result = 16'd250
         973      :	result = 16'd250
         974      :	result = 16'd250
         975      :	result = 16'd250
         976      :	result = 16'd250
         977      :	result = 16'd250
         978      :	result = 16'd250
         979      :	result = 16'd250
         980      :	result = 16'd250
         981      :	result = 16'd250
         982      :	result = 16'd250
         983      :	result = 16'd250
         984      :	result = 16'd250
         985      :	result = 16'd250
         986      :	result = 16'd250
         987      :	result = 16'd250
         988      :	result = 16'd250
         989      :	result = 16'd250
         990      :	result = 16'd250
         991      :	result = 16'd250
         992      :	result = 16'd250
         993      :	result = 16'd250
         994      :	result = 16'd250
         995      :	result = 16'd250
         996      :	result = 16'd250
         997      :	result = 16'd250
         998      :	result = 16'd250
         999      :	result = 16'd250
         1000     :	result = 16'd250
         1001     :	result = 16'd250
         1002     :	result = 16'd251
         1003     :	result = 16'd251
         1004     :	result = 16'd251
         1005     :	result = 16'd251
         1006     :	result = 16'd251
         1007     :	result = 16'd251
         1008     :	result = 16'd251
         1009     :	result = 16'd251
         1010     :	result = 16'd251
         1011     :	result = 16'd251
         1012     :	result = 16'd251
         1013     :	result = 16'd251
         1014     :	result = 16'd251
         1015     :	result = 16'd251
         1016     :	result = 16'd251
         1017     :	result = 16'd251
         1018     :	result = 16'd251
         1019     :	result = 16'd251
         1020     :	result = 16'd251
         1021     :	result = 16'd251
         1022     :	result = 16'd251
         1023     :	result = 16'd251
         1024     :	result = 16'd251
         1025     :	result = 16'd251
         1026     :	result = 16'd251
         1027     :	result = 16'd251
         1028     :	result = 16'd251
         1029     :	result = 16'd251
         1030     :	result = 16'd251
         1031     :	result = 16'd251
         1032     :	result = 16'd251
         1033     :	result = 16'd251
         1034     :	result = 16'd251
         1035     :	result = 16'd251
         1036     :	result = 16'd251
         1037     :	result = 16'd251
         1038     :	result = 16'd251
         1039     :	result = 16'd251
         1040     :	result = 16'd251
         1041     :	result = 16'd251
         1042     :	result = 16'd251
         1043     :	result = 16'd251
         1044     :	result = 16'd251
         1045     :	result = 16'd251
         1046     :	result = 16'd251
         1047     :	result = 16'd251
         1048     :	result = 16'd251
         1049     :	result = 16'd251
         1050     :	result = 16'd251
         1051     :	result = 16'd251
         1052     :	result = 16'd251
         1053     :	result = 16'd251
         1054     :	result = 16'd251
         1055     :	result = 16'd251
         1056     :	result = 16'd251
         1057     :	result = 16'd251
         1058     :	result = 16'd251
         1059     :	result = 16'd251
         1060     :	result = 16'd252
         1061     :	result = 16'd252
         1062     :	result = 16'd252
         1063     :	result = 16'd252
         1064     :	result = 16'd252
         1065     :	result = 16'd252
         1066     :	result = 16'd252
         1067     :	result = 16'd252
         1068     :	result = 16'd252
         1069     :	result = 16'd252
         1070     :	result = 16'd252
         1071     :	result = 16'd252
         1072     :	result = 16'd252
         1073     :	result = 16'd252
         1074     :	result = 16'd252
         1075     :	result = 16'd252
         1076     :	result = 16'd252
         1077     :	result = 16'd252
         1078     :	result = 16'd252
         1079     :	result = 16'd252
         1080     :	result = 16'd252
         1081     :	result = 16'd252
         1082     :	result = 16'd252
         1083     :	result = 16'd252
         1084     :	result = 16'd252
         1085     :	result = 16'd252
         1086     :	result = 16'd252
         1087     :	result = 16'd252
         1088     :	result = 16'd252
         1089     :	result = 16'd252
         1090     :	result = 16'd252
         1091     :	result = 16'd252
         1092     :	result = 16'd252
         1093     :	result = 16'd252
         1094     :	result = 16'd252
         1095     :	result = 16'd252
         1096     :	result = 16'd252
         1097     :	result = 16'd252
         1098     :	result = 16'd252
         1099     :	result = 16'd252
         1100     :	result = 16'd252
         1101     :	result = 16'd252
         1102     :	result = 16'd252
         1103     :	result = 16'd252
         1104     :	result = 16'd252
         1105     :	result = 16'd252
         1106     :	result = 16'd252
         1107     :	result = 16'd252
         1108     :	result = 16'd252
         1109     :	result = 16'd252
         1110     :	result = 16'd252
         1111     :	result = 16'd252
         1112     :	result = 16'd252
         1113     :	result = 16'd252
         1114     :	result = 16'd252
         1115     :	result = 16'd252
         1116     :	result = 16'd252
         1117     :	result = 16'd252
         1118     :	result = 16'd252
         1119     :	result = 16'd252
         1120     :	result = 16'd252
         1121     :	result = 16'd252
         1122     :	result = 16'd252
         1123     :	result = 16'd252
         1124     :	result = 16'd252
         1125     :	result = 16'd252
         1126     :	result = 16'd252
         1127     :	result = 16'd252
         1128     :	result = 16'd252
         1129     :	result = 16'd252
         1130     :	result = 16'd252
         1131     :	result = 16'd252
         1132     :	result = 16'd252
         1133     :	result = 16'd252
         1134     :	result = 16'd252
         1135     :	result = 16'd253
         1136     :	result = 16'd253
         1137     :	result = 16'd253
         1138     :	result = 16'd253
         1139     :	result = 16'd253
         1140     :	result = 16'd253
         1141     :	result = 16'd253
         1142     :	result = 16'd253
         1143     :	result = 16'd253
         1144     :	result = 16'd253
         1145     :	result = 16'd253
         1146     :	result = 16'd253
         1147     :	result = 16'd253
         1148     :	result = 16'd253
         1149     :	result = 16'd253
         1150     :	result = 16'd253
         1151     :	result = 16'd253
         1152     :	result = 16'd253
         1153     :	result = 16'd253
         1154     :	result = 16'd253
         1155     :	result = 16'd253
         1156     :	result = 16'd253
         1157     :	result = 16'd253
         1158     :	result = 16'd253
         1159     :	result = 16'd253
         1160     :	result = 16'd253
         1161     :	result = 16'd253
         1162     :	result = 16'd253
         1163     :	result = 16'd253
         1164     :	result = 16'd253
         1165     :	result = 16'd253
         1166     :	result = 16'd253
         1167     :	result = 16'd253
         1168     :	result = 16'd253
         1169     :	result = 16'd253
         1170     :	result = 16'd253
         1171     :	result = 16'd253
         1172     :	result = 16'd253
         1173     :	result = 16'd253
         1174     :	result = 16'd253
         1175     :	result = 16'd253
         1176     :	result = 16'd253
         1177     :	result = 16'd253
         1178     :	result = 16'd253
         1179     :	result = 16'd253
         1180     :	result = 16'd253
         1181     :	result = 16'd253
         1182     :	result = 16'd253
         1183     :	result = 16'd253
         1184     :	result = 16'd253
         1185     :	result = 16'd253
         1186     :	result = 16'd253
         1187     :	result = 16'd253
         1188     :	result = 16'd253
         1189     :	result = 16'd253
         1190     :	result = 16'd253
         1191     :	result = 16'd253
         1192     :	result = 16'd253
         1193     :	result = 16'd253
         1194     :	result = 16'd253
         1195     :	result = 16'd253
         1196     :	result = 16'd253
         1197     :	result = 16'd253
         1198     :	result = 16'd253
         1199     :	result = 16'd253
         1200     :	result = 16'd253
         1201     :	result = 16'd253
         1202     :	result = 16'd253
         1203     :	result = 16'd253
         1204     :	result = 16'd253
         1205     :	result = 16'd253
         1206     :	result = 16'd253
         1207     :	result = 16'd253
         1208     :	result = 16'd253
         1209     :	result = 16'd253
         1210     :	result = 16'd253
         1211     :	result = 16'd253
         1212     :	result = 16'd253
         1213     :	result = 16'd253
         1214     :	result = 16'd253
         1215     :	result = 16'd253
         1216     :	result = 16'd253
         1217     :	result = 16'd253
         1218     :	result = 16'd253
         1219     :	result = 16'd253
         1220     :	result = 16'd253
         1221     :	result = 16'd253
         1222     :	result = 16'd253
         1223     :	result = 16'd253
         1224     :	result = 16'd253
         1225     :	result = 16'd253
         1226     :	result = 16'd253
         1227     :	result = 16'd253
         1228     :	result = 16'd253
         1229     :	result = 16'd253
         1230     :	result = 16'd253
         1231     :	result = 16'd253
         1232     :	result = 16'd253
         1233     :	result = 16'd253
         1234     :	result = 16'd253
         1235     :	result = 16'd253
         1236     :	result = 16'd253
         1237     :	result = 16'd253
         1238     :	result = 16'd253
         1239     :	result = 16'd253
         1240     :	result = 16'd254
         1241     :	result = 16'd254
         1242     :	result = 16'd254
         1243     :	result = 16'd254
         1244     :	result = 16'd254
         1245     :	result = 16'd254
         1246     :	result = 16'd254
         1247     :	result = 16'd254
         1248     :	result = 16'd254
         1249     :	result = 16'd254
         1250     :	result = 16'd254
         1251     :	result = 16'd254
         1252     :	result = 16'd254
         1253     :	result = 16'd254
         1254     :	result = 16'd254
         1255     :	result = 16'd254
         1256     :	result = 16'd254
         1257     :	result = 16'd254
         1258     :	result = 16'd254
         1259     :	result = 16'd254
         1260     :	result = 16'd254
         1261     :	result = 16'd254
         1262     :	result = 16'd254
         1263     :	result = 16'd254
         1264     :	result = 16'd254
         1265     :	result = 16'd254
         1266     :	result = 16'd254
         1267     :	result = 16'd254
         1268     :	result = 16'd254
         1269     :	result = 16'd254
         1270     :	result = 16'd254
         1271     :	result = 16'd254
         1272     :	result = 16'd254
         1273     :	result = 16'd254
         1274     :	result = 16'd254
         1275     :	result = 16'd254
         1276     :	result = 16'd254
         1277     :	result = 16'd254
         1278     :	result = 16'd254
         1279     :	result = 16'd254
         1280     :	result = 16'd254
         1281     :	result = 16'd254
         1282     :	result = 16'd254
         1283     :	result = 16'd254
         1284     :	result = 16'd254
         1285     :	result = 16'd254
         1286     :	result = 16'd254
         1287     :	result = 16'd254
         1288     :	result = 16'd254
         1289     :	result = 16'd254
         1290     :	result = 16'd254
         1291     :	result = 16'd254
         1292     :	result = 16'd254
         1293     :	result = 16'd254
         1294     :	result = 16'd254
         1295     :	result = 16'd254
         1296     :	result = 16'd254
         1297     :	result = 16'd254
         1298     :	result = 16'd254
         1299     :	result = 16'd254
         1300     :	result = 16'd254
         1301     :	result = 16'd254
         1302     :	result = 16'd254
         1303     :	result = 16'd254
         1304     :	result = 16'd254
         1305     :	result = 16'd254
         1306     :	result = 16'd254
         1307     :	result = 16'd254
         1308     :	result = 16'd254
         1309     :	result = 16'd254
         1310     :	result = 16'd254
         1311     :	result = 16'd254
         1312     :	result = 16'd254
         1313     :	result = 16'd254
         1314     :	result = 16'd254
         1315     :	result = 16'd254
         1316     :	result = 16'd254
         1317     :	result = 16'd254
         1318     :	result = 16'd254
         1319     :	result = 16'd254
         1320     :	result = 16'd254
         1321     :	result = 16'd254
         1322     :	result = 16'd254
         1323     :	result = 16'd254
         1324     :	result = 16'd254
         1325     :	result = 16'd254
         1326     :	result = 16'd254
         1327     :	result = 16'd254
         1328     :	result = 16'd254
         1329     :	result = 16'd254
         1330     :	result = 16'd254
         1331     :	result = 16'd254
         1332     :	result = 16'd254
         1333     :	result = 16'd254
         1334     :	result = 16'd254
         1335     :	result = 16'd254
         1336     :	result = 16'd254
         1337     :	result = 16'd254
         1338     :	result = 16'd254
         1339     :	result = 16'd254
         1340     :	result = 16'd254
         1341     :	result = 16'd254
         1342     :	result = 16'd254
         1343     :	result = 16'd254
         1344     :	result = 16'd254
         1345     :	result = 16'd254
         1346     :	result = 16'd254
         1347     :	result = 16'd254
         1348     :	result = 16'd254
         1349     :	result = 16'd254
         1350     :	result = 16'd254
         1351     :	result = 16'd254
         1352     :	result = 16'd254
         1353     :	result = 16'd254
         1354     :	result = 16'd254
         1355     :	result = 16'd254
         1356     :	result = 16'd254
         1357     :	result = 16'd254
         1358     :	result = 16'd254
         1359     :	result = 16'd254
         1360     :	result = 16'd254
         1361     :	result = 16'd254
         1362     :	result = 16'd254
         1363     :	result = 16'd254
         1364     :	result = 16'd254
         1365     :	result = 16'd254
         1366     :	result = 16'd254
         1367     :	result = 16'd254
         1368     :	result = 16'd254
         1369     :	result = 16'd254
         1370     :	result = 16'd254
         1371     :	result = 16'd254
         1372     :	result = 16'd254
         1373     :	result = 16'd254
         1374     :	result = 16'd254
         1375     :	result = 16'd254
         1376     :	result = 16'd254
         1377     :	result = 16'd254
         1378     :	result = 16'd254
         1379     :	result = 16'd254
         1380     :	result = 16'd254
         1381     :	result = 16'd254
         1382     :	result = 16'd254
         1383     :	result = 16'd254
         1384     :	result = 16'd254
         1385     :	result = 16'd254
         1386     :	result = 16'd254
         1387     :	result = 16'd254
         1388     :	result = 16'd254
         1389     :	result = 16'd254
         1390     :	result = 16'd254
         1391     :	result = 16'd254
         1392     :	result = 16'd254
         1393     :	result = 16'd254
         1394     :	result = 16'd254
         1395     :	result = 16'd254
         1396     :	result = 16'd254
         1397     :	result = 16'd254
         1398     :	result = 16'd254
         1399     :	result = 16'd254
         1400     :	result = 16'd254
         1401     :	result = 16'd254
         1402     :	result = 16'd254
         1403     :	result = 16'd254
         1404     :	result = 16'd254
         1405     :	result = 16'd254
         1406     :	result = 16'd254
         1407     :	result = 16'd254
         1408     :	result = 16'd254
         1409     :	result = 16'd254
         1410     :	result = 16'd254
         1411     :	result = 16'd254
         1412     :	result = 16'd254
         1413     :	result = 16'd254
         1414     :	result = 16'd254
         1415     :	result = 16'd254
         1416     :	result = 16'd254
         1417     :	result = 16'd254
         1418     :	result = 16'd255
         1419     :	result = 16'd255
         1420     :	result = 16'd255
         1421     :	result = 16'd255
         1422     :	result = 16'd255
         1423     :	result = 16'd255
         1424     :	result = 16'd255
         1425     :	result = 16'd255
         1426     :	result = 16'd255
         1427     :	result = 16'd255
         1428     :	result = 16'd255
         1429     :	result = 16'd255
         1430     :	result = 16'd255
         1431     :	result = 16'd255
         1432     :	result = 16'd255
         1433     :	result = 16'd255
         1434     :	result = 16'd255
         1435     :	result = 16'd255
         1436     :	result = 16'd255
         1437     :	result = 16'd255
         1438     :	result = 16'd255
         1439     :	result = 16'd255
         1440     :	result = 16'd255
         1441     :	result = 16'd255
         1442     :	result = 16'd255
         1443     :	result = 16'd255
         1444     :	result = 16'd255
         1445     :	result = 16'd255
         1446     :	result = 16'd255
         1447     :	result = 16'd255
         1448     :	result = 16'd255
         1449     :	result = 16'd255
         1450     :	result = 16'd255
         1451     :	result = 16'd255
         1452     :	result = 16'd255
         1453     :	result = 16'd255
         1454     :	result = 16'd255
         1455     :	result = 16'd255
         1456     :	result = 16'd255
         1457     :	result = 16'd255
         1458     :	result = 16'd255
         1459     :	result = 16'd255
         1460     :	result = 16'd255
         1461     :	result = 16'd255
         1462     :	result = 16'd255
         1463     :	result = 16'd255
         1464     :	result = 16'd255
         1465     :	result = 16'd255
         1466     :	result = 16'd255
         1467     :	result = 16'd255
         1468     :	result = 16'd255
         1469     :	result = 16'd255
         1470     :	result = 16'd255
         1471     :	result = 16'd255
         1472     :	result = 16'd255
         1473     :	result = 16'd255
         1474     :	result = 16'd255
         1475     :	result = 16'd255
         1476     :	result = 16'd255
         1477     :	result = 16'd255
         1478     :	result = 16'd255
         1479     :	result = 16'd255
         1480     :	result = 16'd255
         1481     :	result = 16'd255
         1482     :	result = 16'd255
         1483     :	result = 16'd255
         1484     :	result = 16'd255
         1485     :	result = 16'd255
         1486     :	result = 16'd255
         1487     :	result = 16'd255
         1488     :	result = 16'd255
         1489     :	result = 16'd255
         1490     :	result = 16'd255
         1491     :	result = 16'd255
         1492     :	result = 16'd255
         1493     :	result = 16'd255
         1494     :	result = 16'd255
         1495     :	result = 16'd255
         1496     :	result = 16'd255
         1497     :	result = 16'd255
         1498     :	result = 16'd255
         1499     :	result = 16'd255
         1500     :	result = 16'd255
         1501     :	result = 16'd255
         1502     :	result = 16'd255
         1503     :	result = 16'd255
         1504     :	result = 16'd255
         1505     :	result = 16'd255
         1506     :	result = 16'd255
         1507     :	result = 16'd255
         1508     :	result = 16'd255
         1509     :	result = 16'd255
         1510     :	result = 16'd255
         1511     :	result = 16'd255
         1512     :	result = 16'd255
         1513     :	result = 16'd255
         1514     :	result = 16'd255
         1515     :	result = 16'd255
         1516     :	result = 16'd255
         1517     :	result = 16'd255
         1518     :	result = 16'd255
         1519     :	result = 16'd255
         1520     :	result = 16'd255
         1521     :	result = 16'd255
         1522     :	result = 16'd255
         1523     :	result = 16'd255
         1524     :	result = 16'd255
         1525     :	result = 16'd255
         1526     :	result = 16'd255
         1527     :	result = 16'd255
         1528     :	result = 16'd255
         1529     :	result = 16'd255
         1530     :	result = 16'd255
         1531     :	result = 16'd255
         1532     :	result = 16'd255
         1533     :	result = 16'd255
         1534     :	result = 16'd255
         1535     :	result = 16'd255
         1536     :	result = 16'd255
         1537     :	result = 16'd255
         1538     :	result = 16'd255
         1539     :	result = 16'd255
         1540     :	result = 16'd255
         1541     :	result = 16'd255
         1542     :	result = 16'd255
         1543     :	result = 16'd255
         1544     :	result = 16'd255
         1545     :	result = 16'd255
         1546     :	result = 16'd255
         1547     :	result = 16'd255
         1548     :	result = 16'd255
         1549     :	result = 16'd255
         1550     :	result = 16'd255
         1551     :	result = 16'd255
         1552     :	result = 16'd255
         1553     :	result = 16'd255
         1554     :	result = 16'd255
         1555     :	result = 16'd255
         1556     :	result = 16'd255
         1557     :	result = 16'd255
         1558     :	result = 16'd255
         1559     :	result = 16'd255
         1560     :	result = 16'd255
         1561     :	result = 16'd255
         1562     :	result = 16'd255
         1563     :	result = 16'd255
         1564     :	result = 16'd255
         1565     :	result = 16'd255
         1566     :	result = 16'd255
         1567     :	result = 16'd255
         1568     :	result = 16'd255
         1569     :	result = 16'd255
         1570     :	result = 16'd255
         1571     :	result = 16'd255
         1572     :	result = 16'd255
         1573     :	result = 16'd255
         1574     :	result = 16'd255
         1575     :	result = 16'd255
         1576     :	result = 16'd255
         1577     :	result = 16'd255
         1578     :	result = 16'd255
         1579     :	result = 16'd255
         1580     :	result = 16'd255
         1581     :	result = 16'd255
         1582     :	result = 16'd255
         1583     :	result = 16'd255
         1584     :	result = 16'd255
         1585     :	result = 16'd255
         1586     :	result = 16'd255
         1587     :	result = 16'd255
         1588     :	result = 16'd255
         1589     :	result = 16'd255
         1590     :	result = 16'd255
         1591     :	result = 16'd255
         1592     :	result = 16'd255
         1593     :	result = 16'd255
         1594     :	result = 16'd255
         1595     :	result = 16'd255
         1596     :	result = 16'd255
         1597     :	result = 16'd255
         1598     :	result = 16'd255
         1599     :	result = 16'd255
         1600     :	result = 16'd255
         1601     :	result = 16'd255
         1602     :	result = 16'd255
         1603     :	result = 16'd255
         1604     :	result = 16'd255
         1605     :	result = 16'd255
         1606     :	result = 16'd255
         1607     :	result = 16'd255
         1608     :	result = 16'd255
         1609     :	result = 16'd255
         1610     :	result = 16'd255
         1611     :	result = 16'd255
         1612     :	result = 16'd255
         1613     :	result = 16'd255
         1614     :	result = 16'd255
         1615     :	result = 16'd255
         1616     :	result = 16'd255
         1617     :	result = 16'd255
         1618     :	result = 16'd255
         1619     :	result = 16'd255
         1620     :	result = 16'd255
         1621     :	result = 16'd255
         1622     :	result = 16'd255
         1623     :	result = 16'd255
         1624     :	result = 16'd255
         1625     :	result = 16'd255
         1626     :	result = 16'd255
         1627     :	result = 16'd255
         1628     :	result = 16'd255
         1629     :	result = 16'd255
         1630     :	result = 16'd255
         1631     :	result = 16'd255
         1632     :	result = 16'd255
         1633     :	result = 16'd255
         1634     :	result = 16'd255
         1635     :	result = 16'd255
         1636     :	result = 16'd255
         1637     :	result = 16'd255
         1638     :	result = 16'd255
         1639     :	result = 16'd255
         1640     :	result = 16'd255
         1641     :	result = 16'd255
         1642     :	result = 16'd255
         1643     :	result = 16'd255
         1644     :	result = 16'd255
         1645     :	result = 16'd255
         1646     :	result = 16'd255
         1647     :	result = 16'd255
         1648     :	result = 16'd255
         1649     :	result = 16'd255
         1650     :	result = 16'd255
         1651     :	result = 16'd255
         1652     :	result = 16'd255
         1653     :	result = 16'd255
         1654     :	result = 16'd255
         1655     :	result = 16'd255
         1656     :	result = 16'd255
         1657     :	result = 16'd255
         1658     :	result = 16'd255
         1659     :	result = 16'd255
         1660     :	result = 16'd255
         1661     :	result = 16'd255
         1662     :	result = 16'd255
         1663     :	result = 16'd255
         1664     :	result = 16'd255
         1665     :	result = 16'd255
         1666     :	result = 16'd255
         1667     :	result = 16'd255
         1668     :	result = 16'd255
         1669     :	result = 16'd255
         1670     :	result = 16'd255
         1671     :	result = 16'd255
         1672     :	result = 16'd255
         1673     :	result = 16'd255
         1674     :	result = 16'd255
         1675     :	result = 16'd255
         1676     :	result = 16'd255
         1677     :	result = 16'd255
         1678     :	result = 16'd255
         1679     :	result = 16'd255
         1680     :	result = 16'd255
         1681     :	result = 16'd255
         1682     :	result = 16'd255
         1683     :	result = 16'd255
         1684     :	result = 16'd255
         1685     :	result = 16'd255
         1686     :	result = 16'd255
         1687     :	result = 16'd255
         1688     :	result = 16'd255
         1689     :	result = 16'd255
         1690     :	result = 16'd255
         1691     :	result = 16'd255
         1692     :	result = 16'd255
         1693     :	result = 16'd255
         1694     :	result = 16'd255
         1695     :	result = 16'd255
         1696     :	result = 16'd255
         1697     :	result = 16'd255
         1698     :	result = 16'd255
         1699     :	result = 16'd255
         1700     :	result = 16'd255
         1701     :	result = 16'd255
         1702     :	result = 16'd255
         1703     :	result = 16'd255
         1704     :	result = 16'd255
         1705     :	result = 16'd255
         1706     :	result = 16'd255
         1707     :	result = 16'd255
         1708     :	result = 16'd255
         1709     :	result = 16'd255
         1710     :	result = 16'd255
         1711     :	result = 16'd255
         1712     :	result = 16'd255
         1713     :	result = 16'd255
         1714     :	result = 16'd255
         1715     :	result = 16'd255
         1716     :	result = 16'd255
         1717     :	result = 16'd255
         1718     :	result = 16'd255
         1719     :	result = 16'd255
         1720     :	result = 16'd255
         1721     :	result = 16'd255
         1722     :	result = 16'd255
         1723     :	result = 16'd255
         1724     :	result = 16'd255
         1725     :	result = 16'd255
         1726     :	result = 16'd255
         1727     :	result = 16'd255
         1728     :	result = 16'd255
         1729     :	result = 16'd255
         1730     :	result = 16'd255
         1731     :	result = 16'd255
         1732     :	result = 16'd255
         1733     :	result = 16'd255
         1734     :	result = 16'd255
         1735     :	result = 16'd255
         1736     :	result = 16'd255
         1737     :	result = 16'd255
         1738     :	result = 16'd255
         1739     :	result = 16'd255
         1740     :	result = 16'd255
         1741     :	result = 16'd255
         1742     :	result = 16'd255
         1743     :	result = 16'd255
         1744     :	result = 16'd255
         1745     :	result = 16'd255
         1746     :	result = 16'd255
         1747     :	result = 16'd255
         1748     :	result = 16'd255
         1749     :	result = 16'd255
         1750     :	result = 16'd255
         1751     :	result = 16'd255
         1752     :	result = 16'd255
         1753     :	result = 16'd255
         1754     :	result = 16'd255
         1755     :	result = 16'd255
         1756     :	result = 16'd255
         1757     :	result = 16'd255
         1758     :	result = 16'd255
         1759     :	result = 16'd255
         1760     :	result = 16'd255
         1761     :	result = 16'd255
         1762     :	result = 16'd255
         1763     :	result = 16'd255
         1764     :	result = 16'd255
         1765     :	result = 16'd255
         1766     :	result = 16'd255
         1767     :	result = 16'd255
         1768     :	result = 16'd255
         1769     :	result = 16'd255
         1770     :	result = 16'd255
         1771     :	result = 16'd255
         1772     :	result = 16'd255
         1773     :	result = 16'd255
         1774     :	result = 16'd255
         1775     :	result = 16'd255
         1776     :	result = 16'd255
         1777     :	result = 16'd255
         1778     :	result = 16'd255
         1779     :	result = 16'd255
         1780     :	result = 16'd255
         1781     :	result = 16'd255
         1782     :	result = 16'd255
         1783     :	result = 16'd255
         1784     :	result = 16'd255
         1785     :	result = 16'd255
         1786     :	result = 16'd255
         1787     :	result = 16'd255
         1788     :	result = 16'd255
         1789     :	result = 16'd255
         1790     :	result = 16'd255
         1791     :	result = 16'd255

      endcase
   end

>>>>>>> 60c253bde832c92c80c6fb67bf56cd0ecd0211f4
endmodule