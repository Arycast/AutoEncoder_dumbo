//////////////////////////////////////////////////////////////////////////////////
// Engineer    : Achmad novel, Fauzan Ibrahim, Nicholas Teffandi
// Design Name : Autoencoder
// Module Name : sigmoid_diff_lut
// Project Name: Autoencoder
//////////////////////////////////////////////////////////////////////////////////

// Input and Output is Unsigned

module sigmoid_diff_lut (
   input wire [15:0] addr,
   output reg [15:0] result
);

   always @(*) begin
      
      case (addr)
         63744    :	result = 16'd0;
         63745    :	result = 16'd0;
         63746    :	result = 16'd0;
         63747    :	result = 16'd0;
         63748    :	result = 16'd0;
         63749    :	result = 16'd0;
         63750    :	result = 16'd0;
         63751    :	result = 16'd0;
         63752    :	result = 16'd0;
         63753    :	result = 16'd0;
         63754    :	result = 16'd0;
         63755    :	result = 16'd0;
         63756    :	result = 16'd0;
         63757    :	result = 16'd0;
         63758    :	result = 16'd0;
         63759    :	result = 16'd0;
         63760    :	result = 16'd0;
         63761    :	result = 16'd0;
         63762    :	result = 16'd0;
         63763    :	result = 16'd0;
         63764    :	result = 16'd0;
         63765    :	result = 16'd0;
         63766    :	result = 16'd0;
         63767    :	result = 16'd0;
         63768    :	result = 16'd0;
         63769    :	result = 16'd0;
         63770    :	result = 16'd0;
         63771    :	result = 16'd0;
         63772    :	result = 16'd0;
         63773    :	result = 16'd0;
         63774    :	result = 16'd0;
         63775    :	result = 16'd0;
         63776    :	result = 16'd0;
         63777    :	result = 16'd0;
         63778    :	result = 16'd0;
         63779    :	result = 16'd0;
         63780    :	result = 16'd0;
         63781    :	result = 16'd0;
         63782    :	result = 16'd0;
         63783    :	result = 16'd0;
         63784    :	result = 16'd0;
         63785    :	result = 16'd0;
         63786    :	result = 16'd0;
         63787    :	result = 16'd0;
         63788    :	result = 16'd0;
         63789    :	result = 16'd0;
         63790    :	result = 16'd0;
         63791    :	result = 16'd0;
         63792    :	result = 16'd0;
         63793    :	result = 16'd0;
         63794    :	result = 16'd0;
         63795    :	result = 16'd0;
         63796    :	result = 16'd0;
         63797    :	result = 16'd0;
         63798    :	result = 16'd0;
         63799    :	result = 16'd0;
         63800    :	result = 16'd0;
         63801    :	result = 16'd0;
         63802    :	result = 16'd0;
         63803    :	result = 16'd0;
         63804    :	result = 16'd0;
         63805    :	result = 16'd0;
         63806    :	result = 16'd0;
         63807    :	result = 16'd0;
         63808    :	result = 16'd0;
         63809    :	result = 16'd0;
         63810    :	result = 16'd0;
         63811    :	result = 16'd0;
         63812    :	result = 16'd0;
         63813    :	result = 16'd0;
         63814    :	result = 16'd0;
         63815    :	result = 16'd0;
         63816    :	result = 16'd0;
         63817    :	result = 16'd0;
         63818    :	result = 16'd0;
         63819    :	result = 16'd0;
         63820    :	result = 16'd0;
         63821    :	result = 16'd0;
         63822    :	result = 16'd0;
         63823    :	result = 16'd0;
         63824    :	result = 16'd0;
         63825    :	result = 16'd0;
         63826    :	result = 16'd0;
         63827    :	result = 16'd0;
         63828    :	result = 16'd0;
         63829    :	result = 16'd0;
         63830    :	result = 16'd0;
         63831    :	result = 16'd0;
         63832    :	result = 16'd0;
         63833    :	result = 16'd0;
         63834    :	result = 16'd0;
         63835    :	result = 16'd0;
         63836    :	result = 16'd0;
         63837    :	result = 16'd0;
         63838    :	result = 16'd0;
         63839    :	result = 16'd0;
         63840    :	result = 16'd0;
         63841    :	result = 16'd0;
         63842    :	result = 16'd0;
         63843    :	result = 16'd0;
         63844    :	result = 16'd0;
         63845    :	result = 16'd0;
         63846    :	result = 16'd0;
         63847    :	result = 16'd0;
         63848    :	result = 16'd0;
         63849    :	result = 16'd0;
         63850    :	result = 16'd0;
         63851    :	result = 16'd0;
         63852    :	result = 16'd0;
         63853    :	result = 16'd0;
         63854    :	result = 16'd0;
         63855    :	result = 16'd0;
         63856    :	result = 16'd0;
         63857    :	result = 16'd0;
         63858    :	result = 16'd0;
         63859    :	result = 16'd0;
         63860    :	result = 16'd0;
         63861    :	result = 16'd0;
         63862    :	result = 16'd0;
         63863    :	result = 16'd0;
         63864    :	result = 16'd0;
         63865    :	result = 16'd0;
         63866    :	result = 16'd0;
         63867    :	result = 16'd0;
         63868    :	result = 16'd0;
         63869    :	result = 16'd0;
         63870    :	result = 16'd0;
         63871    :	result = 16'd0;
         63872    :	result = 16'd0;
         63873    :	result = 16'd0;
         63874    :	result = 16'd0;
         63875    :	result = 16'd0;
         63876    :	result = 16'd0;
         63877    :	result = 16'd0;
         63878    :	result = 16'd0;
         63879    :	result = 16'd0;
         63880    :	result = 16'd0;
         63881    :	result = 16'd0;
         63882    :	result = 16'd0;
         63883    :	result = 16'd0;
         63884    :	result = 16'd0;
         63885    :	result = 16'd0;
         63886    :	result = 16'd0;
         63887    :	result = 16'd0;
         63888    :	result = 16'd0;
         63889    :	result = 16'd0;
         63890    :	result = 16'd0;
         63891    :	result = 16'd0;
         63892    :	result = 16'd0;
         63893    :	result = 16'd0;
         63894    :	result = 16'd0;
         63895    :	result = 16'd0;
         63896    :	result = 16'd0;
         63897    :	result = 16'd0;
         63898    :	result = 16'd0;
         63899    :	result = 16'd0;
         63900    :	result = 16'd0;
         63901    :	result = 16'd0;
         63902    :	result = 16'd0;
         63903    :	result = 16'd0;
         63904    :	result = 16'd0;
         63905    :	result = 16'd0;
         63906    :	result = 16'd0;
         63907    :	result = 16'd0;
         63908    :	result = 16'd0;
         63909    :	result = 16'd0;
         63910    :	result = 16'd0;
         63911    :	result = 16'd0;
         63912    :	result = 16'd0;
         63913    :	result = 16'd0;
         63914    :	result = 16'd0;
         63915    :	result = 16'd0;
         63916    :	result = 16'd0;
         63917    :	result = 16'd0;
         63918    :	result = 16'd0;
         63919    :	result = 16'd0;
         63920    :	result = 16'd0;
         63921    :	result = 16'd0;
         63922    :	result = 16'd0;
         63923    :	result = 16'd0;
         63924    :	result = 16'd0;
         63925    :	result = 16'd0;
         63926    :	result = 16'd0;
         63927    :	result = 16'd0;
         63928    :	result = 16'd0;
         63929    :	result = 16'd0;
         63930    :	result = 16'd0;
         63931    :	result = 16'd0;
         63932    :	result = 16'd0;
         63933    :	result = 16'd0;
         63934    :	result = 16'd0;
         63935    :	result = 16'd0;
         63936    :	result = 16'd0;
         63937    :	result = 16'd0;
         63938    :	result = 16'd0;
         63939    :	result = 16'd0;
         63940    :	result = 16'd0;
         63941    :	result = 16'd0;
         63942    :	result = 16'd0;
         63943    :	result = 16'd0;
         63944    :	result = 16'd0;
         63945    :	result = 16'd0;
         63946    :	result = 16'd0;
         63947    :	result = 16'd0;
         63948    :	result = 16'd0;
         63949    :	result = 16'd0;
         63950    :	result = 16'd0;
         63951    :	result = 16'd0;
         63952    :	result = 16'd0;
         63953    :	result = 16'd0;
         63954    :	result = 16'd0;
         63955    :	result = 16'd0;
         63956    :	result = 16'd0;
         63957    :	result = 16'd0;
         63958    :	result = 16'd0;
         63959    :	result = 16'd0;
         63960    :	result = 16'd0;
         63961    :	result = 16'd0;
         63962    :	result = 16'd0;
         63963    :	result = 16'd0;
         63964    :	result = 16'd0;
         63965    :	result = 16'd0;
         63966    :	result = 16'd0;
         63967    :	result = 16'd0;
         63968    :	result = 16'd0;
         63969    :	result = 16'd0;
         63970    :	result = 16'd0;
         63971    :	result = 16'd0;
         63972    :	result = 16'd0;
         63973    :	result = 16'd0;
         63974    :	result = 16'd0;
         63975    :	result = 16'd0;
         63976    :	result = 16'd0;
         63977    :	result = 16'd0;
         63978    :	result = 16'd0;
         63979    :	result = 16'd0;
         63980    :	result = 16'd0;
         63981    :	result = 16'd0;
         63982    :	result = 16'd0;
         63983    :	result = 16'd0;
         63984    :	result = 16'd0;
         63985    :	result = 16'd0;
         63986    :	result = 16'd0;
         63987    :	result = 16'd0;
         63988    :	result = 16'd0;
         63989    :	result = 16'd0;
         63990    :	result = 16'd0;
         63991    :	result = 16'd0;
         63992    :	result = 16'd0;
         63993    :	result = 16'd0;
         63994    :	result = 16'd0;
         63995    :	result = 16'd0;
         63996    :	result = 16'd0;
         63997    :	result = 16'd0;
         63998    :	result = 16'd0;
         63999    :	result = 16'd0;
         64000    :	result = 16'd0;
         64001    :	result = 16'd0;
         64002    :	result = 16'd0;
         64003    :	result = 16'd0;
         64004    :	result = 16'd0;
         64005    :	result = 16'd0;
         64006    :	result = 16'd0;
         64007    :	result = 16'd0;
         64008    :	result = 16'd0;
         64009    :	result = 16'd0;
         64010    :	result = 16'd0;
         64011    :	result = 16'd0;
         64012    :	result = 16'd0;
         64013    :	result = 16'd0;
         64014    :	result = 16'd0;
         64015    :	result = 16'd0;
         64016    :	result = 16'd0;
         64017    :	result = 16'd0;
         64018    :	result = 16'd0;
         64019    :	result = 16'd0;
         64020    :	result = 16'd0;
         64021    :	result = 16'd0;
         64022    :	result = 16'd0;
         64023    :	result = 16'd0;
         64024    :	result = 16'd0;
         64025    :	result = 16'd0;
         64026    :	result = 16'd0;
         64027    :	result = 16'd0;
         64028    :	result = 16'd0;
         64029    :	result = 16'd0;
         64030    :	result = 16'd0;
         64031    :	result = 16'd0;
         64032    :	result = 16'd0;
         64033    :	result = 16'd0;
         64034    :	result = 16'd0;
         64035    :	result = 16'd0;
         64036    :	result = 16'd0;
         64037    :	result = 16'd0;
         64038    :	result = 16'd0;
         64039    :	result = 16'd0;
         64040    :	result = 16'd0;
         64041    :	result = 16'd0;
         64042    :	result = 16'd0;
         64043    :	result = 16'd0;
         64044    :	result = 16'd0;
         64045    :	result = 16'd0;
         64046    :	result = 16'd0;
         64047    :	result = 16'd0;
         64048    :	result = 16'd0;
         64049    :	result = 16'd0;
         64050    :	result = 16'd0;
         64051    :	result = 16'd0;
         64052    :	result = 16'd0;
         64053    :	result = 16'd0;
         64054    :	result = 16'd0;
         64055    :	result = 16'd0;
         64056    :	result = 16'd0;
         64057    :	result = 16'd0;
         64058    :	result = 16'd0;
         64059    :	result = 16'd0;
         64060    :	result = 16'd0;
         64061    :	result = 16'd0;
         64062    :	result = 16'd0;
         64063    :	result = 16'd0;
         64064    :	result = 16'd0;
         64065    :	result = 16'd0;
         64066    :	result = 16'd0;
         64067    :	result = 16'd0;
         64068    :	result = 16'd0;
         64069    :	result = 16'd0;
         64070    :	result = 16'd0;
         64071    :	result = 16'd0;
         64072    :	result = 16'd0;
         64073    :	result = 16'd0;
         64074    :	result = 16'd0;
         64075    :	result = 16'd0;
         64076    :	result = 16'd0;
         64077    :	result = 16'd0;
         64078    :	result = 16'd0;
         64079    :	result = 16'd0;
         64080    :	result = 16'd0;
         64081    :	result = 16'd0;
         64082    :	result = 16'd0;
         64083    :	result = 16'd0;
         64084    :	result = 16'd0;
         64085    :	result = 16'd0;
         64086    :	result = 16'd0;
         64087    :	result = 16'd0;
         64088    :	result = 16'd0;
         64089    :	result = 16'd0;
         64090    :	result = 16'd0;
         64091    :	result = 16'd0;
         64092    :	result = 16'd0;
         64093    :	result = 16'd0;
         64094    :	result = 16'd0;
         64095    :	result = 16'd0;
         64096    :	result = 16'd0;
         64097    :	result = 16'd0;
         64098    :	result = 16'd0;
         64099    :	result = 16'd0;
         64100    :	result = 16'd0;
         64101    :	result = 16'd0;
         64102    :	result = 16'd0;
         64103    :	result = 16'd0;
         64104    :	result = 16'd0;
         64105    :	result = 16'd0;
         64106    :	result = 16'd0;
         64107    :	result = 16'd0;
         64108    :	result = 16'd0;
         64109    :	result = 16'd0;
         64110    :	result = 16'd0;
         64111    :	result = 16'd0;
         64112    :	result = 16'd0;
         64113    :	result = 16'd0;
         64114    :	result = 16'd0;
         64115    :	result = 16'd0;
         64116    :	result = 16'd0;
         64117    :	result = 16'd0;
         64118    :	result = 16'd1;
         64119    :	result = 16'd1;
         64120    :	result = 16'd1;
         64121    :	result = 16'd1;
         64122    :	result = 16'd1;
         64123    :	result = 16'd1;
         64124    :	result = 16'd1;
         64125    :	result = 16'd1;
         64126    :	result = 16'd1;
         64127    :	result = 16'd1;
         64128    :	result = 16'd1;
         64129    :	result = 16'd1;
         64130    :	result = 16'd1;
         64131    :	result = 16'd1;
         64132    :	result = 16'd1;
         64133    :	result = 16'd1;
         64134    :	result = 16'd1;
         64135    :	result = 16'd1;
         64136    :	result = 16'd1;
         64137    :	result = 16'd1;
         64138    :	result = 16'd1;
         64139    :	result = 16'd1;
         64140    :	result = 16'd1;
         64141    :	result = 16'd1;
         64142    :	result = 16'd1;
         64143    :	result = 16'd1;
         64144    :	result = 16'd1;
         64145    :	result = 16'd1;
         64146    :	result = 16'd1;
         64147    :	result = 16'd1;
         64148    :	result = 16'd1;
         64149    :	result = 16'd1;
         64150    :	result = 16'd1;
         64151    :	result = 16'd1;
         64152    :	result = 16'd1;
         64153    :	result = 16'd1;
         64154    :	result = 16'd1;
         64155    :	result = 16'd1;
         64156    :	result = 16'd1;
         64157    :	result = 16'd1;
         64158    :	result = 16'd1;
         64159    :	result = 16'd1;
         64160    :	result = 16'd1;
         64161    :	result = 16'd1;
         64162    :	result = 16'd1;
         64163    :	result = 16'd1;
         64164    :	result = 16'd1;
         64165    :	result = 16'd1;
         64166    :	result = 16'd1;
         64167    :	result = 16'd1;
         64168    :	result = 16'd1;
         64169    :	result = 16'd1;
         64170    :	result = 16'd1;
         64171    :	result = 16'd1;
         64172    :	result = 16'd1;
         64173    :	result = 16'd1;
         64174    :	result = 16'd1;
         64175    :	result = 16'd1;
         64176    :	result = 16'd1;
         64177    :	result = 16'd1;
         64178    :	result = 16'd1;
         64179    :	result = 16'd1;
         64180    :	result = 16'd1;
         64181    :	result = 16'd1;
         64182    :	result = 16'd1;
         64183    :	result = 16'd1;
         64184    :	result = 16'd1;
         64185    :	result = 16'd1;
         64186    :	result = 16'd1;
         64187    :	result = 16'd1;
         64188    :	result = 16'd1;
         64189    :	result = 16'd1;
         64190    :	result = 16'd1;
         64191    :	result = 16'd1;
         64192    :	result = 16'd1;
         64193    :	result = 16'd1;
         64194    :	result = 16'd1;
         64195    :	result = 16'd1;
         64196    :	result = 16'd1;
         64197    :	result = 16'd1;
         64198    :	result = 16'd1;
         64199    :	result = 16'd1;
         64200    :	result = 16'd1;
         64201    :	result = 16'd1;
         64202    :	result = 16'd1;
         64203    :	result = 16'd1;
         64204    :	result = 16'd1;
         64205    :	result = 16'd1;
         64206    :	result = 16'd1;
         64207    :	result = 16'd1;
         64208    :	result = 16'd1;
         64209    :	result = 16'd1;
         64210    :	result = 16'd1;
         64211    :	result = 16'd1;
         64212    :	result = 16'd1;
         64213    :	result = 16'd1;
         64214    :	result = 16'd1;
         64215    :	result = 16'd1;
         64216    :	result = 16'd1;
         64217    :	result = 16'd1;
         64218    :	result = 16'd1;
         64219    :	result = 16'd1;
         64220    :	result = 16'd1;
         64221    :	result = 16'd1;
         64222    :	result = 16'd1;
         64223    :	result = 16'd1;
         64224    :	result = 16'd1;
         64225    :	result = 16'd1;
         64226    :	result = 16'd1;
         64227    :	result = 16'd1;
         64228    :	result = 16'd1;
         64229    :	result = 16'd1;
         64230    :	result = 16'd1;
         64231    :	result = 16'd1;
         64232    :	result = 16'd1;
         64233    :	result = 16'd1;
         64234    :	result = 16'd1;
         64235    :	result = 16'd1;
         64236    :	result = 16'd1;
         64237    :	result = 16'd1;
         64238    :	result = 16'd1;
         64239    :	result = 16'd1;
         64240    :	result = 16'd1;
         64241    :	result = 16'd1;
         64242    :	result = 16'd1;
         64243    :	result = 16'd1;
         64244    :	result = 16'd1;
         64245    :	result = 16'd1;
         64246    :	result = 16'd1;
         64247    :	result = 16'd1;
         64248    :	result = 16'd1;
         64249    :	result = 16'd1;
         64250    :	result = 16'd1;
         64251    :	result = 16'd1;
         64252    :	result = 16'd1;
         64253    :	result = 16'd1;
         64254    :	result = 16'd1;
         64255    :	result = 16'd1;
         64256    :	result = 16'd1;
         64257    :	result = 16'd1;
         64258    :	result = 16'd1;
         64259    :	result = 16'd1;
         64260    :	result = 16'd1;
         64261    :	result = 16'd1;
         64262    :	result = 16'd1;
         64263    :	result = 16'd1;
         64264    :	result = 16'd1;
         64265    :	result = 16'd1;
         64266    :	result = 16'd1;
         64267    :	result = 16'd1;
         64268    :	result = 16'd1;
         64269    :	result = 16'd1;
         64270    :	result = 16'd1;
         64271    :	result = 16'd1;
         64272    :	result = 16'd1;
         64273    :	result = 16'd1;
         64274    :	result = 16'd1;
         64275    :	result = 16'd1;
         64276    :	result = 16'd1;
         64277    :	result = 16'd1;
         64278    :	result = 16'd1;
         64279    :	result = 16'd1;
         64280    :	result = 16'd1;
         64281    :	result = 16'd1;
         64282    :	result = 16'd1;
         64283    :	result = 16'd1;
         64284    :	result = 16'd1;
         64285    :	result = 16'd1;
         64286    :	result = 16'd1;
         64287    :	result = 16'd1;
         64288    :	result = 16'd1;
         64289    :	result = 16'd1;
         64290    :	result = 16'd1;
         64291    :	result = 16'd1;
         64292    :	result = 16'd1;
         64293    :	result = 16'd1;
         64294    :	result = 16'd1;
         64295    :	result = 16'd1;
         64296    :	result = 16'd1;
         64297    :	result = 16'd2;
         64298    :	result = 16'd2;
         64299    :	result = 16'd2;
         64300    :	result = 16'd2;
         64301    :	result = 16'd2;
         64302    :	result = 16'd2;
         64303    :	result = 16'd2;
         64304    :	result = 16'd2;
         64305    :	result = 16'd2;
         64306    :	result = 16'd2;
         64307    :	result = 16'd2;
         64308    :	result = 16'd2;
         64309    :	result = 16'd2;
         64310    :	result = 16'd2;
         64311    :	result = 16'd2;
         64312    :	result = 16'd2;
         64313    :	result = 16'd2;
         64314    :	result = 16'd2;
         64315    :	result = 16'd2;
         64316    :	result = 16'd2;
         64317    :	result = 16'd2;
         64318    :	result = 16'd2;
         64319    :	result = 16'd2;
         64320    :	result = 16'd2;
         64321    :	result = 16'd2;
         64322    :	result = 16'd2;
         64323    :	result = 16'd2;
         64324    :	result = 16'd2;
         64325    :	result = 16'd2;
         64326    :	result = 16'd2;
         64327    :	result = 16'd2;
         64328    :	result = 16'd2;
         64329    :	result = 16'd2;
         64330    :	result = 16'd2;
         64331    :	result = 16'd2;
         64332    :	result = 16'd2;
         64333    :	result = 16'd2;
         64334    :	result = 16'd2;
         64335    :	result = 16'd2;
         64336    :	result = 16'd2;
         64337    :	result = 16'd2;
         64338    :	result = 16'd2;
         64339    :	result = 16'd2;
         64340    :	result = 16'd2;
         64341    :	result = 16'd2;
         64342    :	result = 16'd2;
         64343    :	result = 16'd2;
         64344    :	result = 16'd2;
         64345    :	result = 16'd2;
         64346    :	result = 16'd2;
         64347    :	result = 16'd2;
         64348    :	result = 16'd2;
         64349    :	result = 16'd2;
         64350    :	result = 16'd2;
         64351    :	result = 16'd2;
         64352    :	result = 16'd2;
         64353    :	result = 16'd2;
         64354    :	result = 16'd2;
         64355    :	result = 16'd2;
         64356    :	result = 16'd2;
         64357    :	result = 16'd2;
         64358    :	result = 16'd2;
         64359    :	result = 16'd2;
         64360    :	result = 16'd2;
         64361    :	result = 16'd2;
         64362    :	result = 16'd2;
         64363    :	result = 16'd2;
         64364    :	result = 16'd2;
         64365    :	result = 16'd2;
         64366    :	result = 16'd2;
         64367    :	result = 16'd2;
         64368    :	result = 16'd2;
         64369    :	result = 16'd2;
         64370    :	result = 16'd2;
         64371    :	result = 16'd2;
         64372    :	result = 16'd2;
         64373    :	result = 16'd2;
         64374    :	result = 16'd2;
         64375    :	result = 16'd2;
         64376    :	result = 16'd2;
         64377    :	result = 16'd2;
         64378    :	result = 16'd2;
         64379    :	result = 16'd2;
         64380    :	result = 16'd2;
         64381    :	result = 16'd2;
         64382    :	result = 16'd2;
         64383    :	result = 16'd2;
         64384    :	result = 16'd2;
         64385    :	result = 16'd2;
         64386    :	result = 16'd2;
         64387    :	result = 16'd2;
         64388    :	result = 16'd2;
         64389    :	result = 16'd2;
         64390    :	result = 16'd2;
         64391    :	result = 16'd2;
         64392    :	result = 16'd2;
         64393    :	result = 16'd2;
         64394    :	result = 16'd2;
         64395    :	result = 16'd2;
         64396    :	result = 16'd2;
         64397    :	result = 16'd2;
         64398    :	result = 16'd2;
         64399    :	result = 16'd2;
         64400    :	result = 16'd2;
         64401    :	result = 16'd2;
         64402    :	result = 16'd2;
         64403    :	result = 16'd3;
         64404    :	result = 16'd3;
         64405    :	result = 16'd3;
         64406    :	result = 16'd3;
         64407    :	result = 16'd3;
         64408    :	result = 16'd3;
         64409    :	result = 16'd3;
         64410    :	result = 16'd3;
         64411    :	result = 16'd3;
         64412    :	result = 16'd3;
         64413    :	result = 16'd3;
         64414    :	result = 16'd3;
         64415    :	result = 16'd3;
         64416    :	result = 16'd3;
         64417    :	result = 16'd3;
         64418    :	result = 16'd3;
         64419    :	result = 16'd3;
         64420    :	result = 16'd3;
         64421    :	result = 16'd3;
         64422    :	result = 16'd3;
         64423    :	result = 16'd3;
         64424    :	result = 16'd3;
         64425    :	result = 16'd3;
         64426    :	result = 16'd3;
         64427    :	result = 16'd3;
         64428    :	result = 16'd3;
         64429    :	result = 16'd3;
         64430    :	result = 16'd3;
         64431    :	result = 16'd3;
         64432    :	result = 16'd3;
         64433    :	result = 16'd3;
         64434    :	result = 16'd3;
         64435    :	result = 16'd3;
         64436    :	result = 16'd3;
         64437    :	result = 16'd3;
         64438    :	result = 16'd3;
         64439    :	result = 16'd3;
         64440    :	result = 16'd3;
         64441    :	result = 16'd3;
         64442    :	result = 16'd3;
         64443    :	result = 16'd3;
         64444    :	result = 16'd3;
         64445    :	result = 16'd3;
         64446    :	result = 16'd3;
         64447    :	result = 16'd3;
         64448    :	result = 16'd3;
         64449    :	result = 16'd3;
         64450    :	result = 16'd3;
         64451    :	result = 16'd3;
         64452    :	result = 16'd3;
         64453    :	result = 16'd3;
         64454    :	result = 16'd3;
         64455    :	result = 16'd3;
         64456    :	result = 16'd3;
         64457    :	result = 16'd3;
         64458    :	result = 16'd3;
         64459    :	result = 16'd3;
         64460    :	result = 16'd3;
         64461    :	result = 16'd3;
         64462    :	result = 16'd3;
         64463    :	result = 16'd3;
         64464    :	result = 16'd3;
         64465    :	result = 16'd3;
         64466    :	result = 16'd3;
         64467    :	result = 16'd3;
         64468    :	result = 16'd3;
         64469    :	result = 16'd3;
         64470    :	result = 16'd3;
         64471    :	result = 16'd3;
         64472    :	result = 16'd3;
         64473    :	result = 16'd3;
         64474    :	result = 16'd3;
         64475    :	result = 16'd3;
         64476    :	result = 16'd3;
         64477    :	result = 16'd3;
         64478    :	result = 16'd3;
         64479    :	result = 16'd4;
         64480    :	result = 16'd4;
         64481    :	result = 16'd4;
         64482    :	result = 16'd4;
         64483    :	result = 16'd4;
         64484    :	result = 16'd4;
         64485    :	result = 16'd4;
         64486    :	result = 16'd4;
         64487    :	result = 16'd4;
         64488    :	result = 16'd4;
         64489    :	result = 16'd4;
         64490    :	result = 16'd4;
         64491    :	result = 16'd4;
         64492    :	result = 16'd4;
         64493    :	result = 16'd4;
         64494    :	result = 16'd4;
         64495    :	result = 16'd4;
         64496    :	result = 16'd4;
         64497    :	result = 16'd4;
         64498    :	result = 16'd4;
         64499    :	result = 16'd4;
         64500    :	result = 16'd4;
         64501    :	result = 16'd4;
         64502    :	result = 16'd4;
         64503    :	result = 16'd4;
         64504    :	result = 16'd4;
         64505    :	result = 16'd4;
         64506    :	result = 16'd4;
         64507    :	result = 16'd4;
         64508    :	result = 16'd4;
         64509    :	result = 16'd4;
         64510    :	result = 16'd4;
         64511    :	result = 16'd4;
         64512    :	result = 16'd4;
         64513    :	result = 16'd4;
         64514    :	result = 16'd4;
         64515    :	result = 16'd4;
         64516    :	result = 16'd4;
         64517    :	result = 16'd4;
         64518    :	result = 16'd4;
         64519    :	result = 16'd4;
         64520    :	result = 16'd4;
         64521    :	result = 16'd4;
         64522    :	result = 16'd4;
         64523    :	result = 16'd4;
         64524    :	result = 16'd4;
         64525    :	result = 16'd4;
         64526    :	result = 16'd4;
         64527    :	result = 16'd4;
         64528    :	result = 16'd4;
         64529    :	result = 16'd4;
         64530    :	result = 16'd4;
         64531    :	result = 16'd4;
         64532    :	result = 16'd4;
         64533    :	result = 16'd4;
         64534    :	result = 16'd4;
         64535    :	result = 16'd4;
         64536    :	result = 16'd4;
         64537    :	result = 16'd4;
         64538    :	result = 16'd5;
         64539    :	result = 16'd5;
         64540    :	result = 16'd5;
         64541    :	result = 16'd5;
         64542    :	result = 16'd5;
         64543    :	result = 16'd5;
         64544    :	result = 16'd5;
         64545    :	result = 16'd5;
         64546    :	result = 16'd5;
         64547    :	result = 16'd5;
         64548    :	result = 16'd5;
         64549    :	result = 16'd5;
         64550    :	result = 16'd5;
         64551    :	result = 16'd5;
         64552    :	result = 16'd5;
         64553    :	result = 16'd5;
         64554    :	result = 16'd5;
         64555    :	result = 16'd5;
         64556    :	result = 16'd5;
         64557    :	result = 16'd5;
         64558    :	result = 16'd5;
         64559    :	result = 16'd5;
         64560    :	result = 16'd5;
         64561    :	result = 16'd5;
         64562    :	result = 16'd5;
         64563    :	result = 16'd5;
         64564    :	result = 16'd5;
         64565    :	result = 16'd5;
         64566    :	result = 16'd5;
         64567    :	result = 16'd5;
         64568    :	result = 16'd5;
         64569    :	result = 16'd5;
         64570    :	result = 16'd5;
         64571    :	result = 16'd5;
         64572    :	result = 16'd5;
         64573    :	result = 16'd5;
         64574    :	result = 16'd5;
         64575    :	result = 16'd5;
         64576    :	result = 16'd5;
         64577    :	result = 16'd5;
         64578    :	result = 16'd5;
         64579    :	result = 16'd5;
         64580    :	result = 16'd5;
         64581    :	result = 16'd5;
         64582    :	result = 16'd5;
         64583    :	result = 16'd5;
         64584    :	result = 16'd5;
         64585    :	result = 16'd5;
         64586    :	result = 16'd5;
         64587    :	result = 16'd6;
         64588    :	result = 16'd6;
         64589    :	result = 16'd6;
         64590    :	result = 16'd6;
         64591    :	result = 16'd6;
         64592    :	result = 16'd6;
         64593    :	result = 16'd6;
         64594    :	result = 16'd6;
         64595    :	result = 16'd6;
         64596    :	result = 16'd6;
         64597    :	result = 16'd6;
         64598    :	result = 16'd6;
         64599    :	result = 16'd6;
         64600    :	result = 16'd6;
         64601    :	result = 16'd6;
         64602    :	result = 16'd6;
         64603    :	result = 16'd6;
         64604    :	result = 16'd6;
         64605    :	result = 16'd6;
         64606    :	result = 16'd6;
         64607    :	result = 16'd6;
         64608    :	result = 16'd6;
         64609    :	result = 16'd6;
         64610    :	result = 16'd6;
         64611    :	result = 16'd6;
         64612    :	result = 16'd6;
         64613    :	result = 16'd6;
         64614    :	result = 16'd6;
         64615    :	result = 16'd6;
         64616    :	result = 16'd6;
         64617    :	result = 16'd6;
         64618    :	result = 16'd6;
         64619    :	result = 16'd6;
         64620    :	result = 16'd6;
         64621    :	result = 16'd6;
         64622    :	result = 16'd6;
         64623    :	result = 16'd6;
         64624    :	result = 16'd6;
         64625    :	result = 16'd6;
         64626    :	result = 16'd6;
         64627    :	result = 16'd6;
         64628    :	result = 16'd6;
         64629    :	result = 16'd7;
         64630    :	result = 16'd7;
         64631    :	result = 16'd7;
         64632    :	result = 16'd7;
         64633    :	result = 16'd7;
         64634    :	result = 16'd7;
         64635    :	result = 16'd7;
         64636    :	result = 16'd7;
         64637    :	result = 16'd7;
         64638    :	result = 16'd7;
         64639    :	result = 16'd7;
         64640    :	result = 16'd7;
         64641    :	result = 16'd7;
         64642    :	result = 16'd7;
         64643    :	result = 16'd7;
         64644    :	result = 16'd7;
         64645    :	result = 16'd7;
         64646    :	result = 16'd7;
         64647    :	result = 16'd7;
         64648    :	result = 16'd7;
         64649    :	result = 16'd7;
         64650    :	result = 16'd7;
         64651    :	result = 16'd7;
         64652    :	result = 16'd7;
         64653    :	result = 16'd7;
         64654    :	result = 16'd7;
         64655    :	result = 16'd7;
         64656    :	result = 16'd7;
         64657    :	result = 16'd7;
         64658    :	result = 16'd7;
         64659    :	result = 16'd7;
         64660    :	result = 16'd7;
         64661    :	result = 16'd7;
         64662    :	result = 16'd7;
         64663    :	result = 16'd7;
         64664    :	result = 16'd7;
         64665    :	result = 16'd8;
         64666    :	result = 16'd8;
         64667    :	result = 16'd8;
         64668    :	result = 16'd8;
         64669    :	result = 16'd8;
         64670    :	result = 16'd8;
         64671    :	result = 16'd8;
         64672    :	result = 16'd8;
         64673    :	result = 16'd8;
         64674    :	result = 16'd8;
         64675    :	result = 16'd8;
         64676    :	result = 16'd8;
         64677    :	result = 16'd8;
         64678    :	result = 16'd8;
         64679    :	result = 16'd8;
         64680    :	result = 16'd8;
         64681    :	result = 16'd8;
         64682    :	result = 16'd8;
         64683    :	result = 16'd8;
         64684    :	result = 16'd8;
         64685    :	result = 16'd8;
         64686    :	result = 16'd8;
         64687    :	result = 16'd8;
         64688    :	result = 16'd8;
         64689    :	result = 16'd8;
         64690    :	result = 16'd8;
         64691    :	result = 16'd8;
         64692    :	result = 16'd8;
         64693    :	result = 16'd8;
         64694    :	result = 16'd8;
         64695    :	result = 16'd8;
         64696    :	result = 16'd8;
         64697    :	result = 16'd9;
         64698    :	result = 16'd9;
         64699    :	result = 16'd9;
         64700    :	result = 16'd9;
         64701    :	result = 16'd9;
         64702    :	result = 16'd9;
         64703    :	result = 16'd9;
         64704    :	result = 16'd9;
         64705    :	result = 16'd9;
         64706    :	result = 16'd9;
         64707    :	result = 16'd9;
         64708    :	result = 16'd9;
         64709    :	result = 16'd9;
         64710    :	result = 16'd9;
         64711    :	result = 16'd9;
         64712    :	result = 16'd9;
         64713    :	result = 16'd9;
         64714    :	result = 16'd9;
         64715    :	result = 16'd9;
         64716    :	result = 16'd9;
         64717    :	result = 16'd9;
         64718    :	result = 16'd9;
         64719    :	result = 16'd9;
         64720    :	result = 16'd9;
         64721    :	result = 16'd9;
         64722    :	result = 16'd9;
         64723    :	result = 16'd9;
         64724    :	result = 16'd9;
         64725    :	result = 16'd9;
         64726    :	result = 16'd9;
         64727    :	result = 16'd10;
         64728    :	result = 16'd10;
         64729    :	result = 16'd10;
         64730    :	result = 16'd10;
         64731    :	result = 16'd10;
         64732    :	result = 16'd10;
         64733    :	result = 16'd10;
         64734    :	result = 16'd10;
         64735    :	result = 16'd10;
         64736    :	result = 16'd10;
         64737    :	result = 16'd10;
         64738    :	result = 16'd10;
         64739    :	result = 16'd10;
         64740    :	result = 16'd10;
         64741    :	result = 16'd10;
         64742    :	result = 16'd10;
         64743    :	result = 16'd10;
         64744    :	result = 16'd10;
         64745    :	result = 16'd10;
         64746    :	result = 16'd10;
         64747    :	result = 16'd10;
         64748    :	result = 16'd10;
         64749    :	result = 16'd10;
         64750    :	result = 16'd10;
         64751    :	result = 16'd10;
         64752    :	result = 16'd10;
         64753    :	result = 16'd11;
         64754    :	result = 16'd11;
         64755    :	result = 16'd11;
         64756    :	result = 16'd11;
         64757    :	result = 16'd11;
         64758    :	result = 16'd11;
         64759    :	result = 16'd11;
         64760    :	result = 16'd11;
         64761    :	result = 16'd11;
         64762    :	result = 16'd11;
         64763    :	result = 16'd11;
         64764    :	result = 16'd11;
         64765    :	result = 16'd11;
         64766    :	result = 16'd11;
         64767    :	result = 16'd11;
         64768    :	result = 16'd11;
         64769    :	result = 16'd11;
         64770    :	result = 16'd11;
         64771    :	result = 16'd11;
         64772    :	result = 16'd11;
         64773    :	result = 16'd11;
         64774    :	result = 16'd11;
         64775    :	result = 16'd11;
         64776    :	result = 16'd11;
         64777    :	result = 16'd11;
         64778    :	result = 16'd12;
         64779    :	result = 16'd12;
         64780    :	result = 16'd12;
         64781    :	result = 16'd12;
         64782    :	result = 16'd12;
         64783    :	result = 16'd12;
         64784    :	result = 16'd12;
         64785    :	result = 16'd12;
         64786    :	result = 16'd12;
         64787    :	result = 16'd12;
         64788    :	result = 16'd12;
         64789    :	result = 16'd12;
         64790    :	result = 16'd12;
         64791    :	result = 16'd12;
         64792    :	result = 16'd12;
         64793    :	result = 16'd12;
         64794    :	result = 16'd12;
         64795    :	result = 16'd12;
         64796    :	result = 16'd12;
         64797    :	result = 16'd12;
         64798    :	result = 16'd12;
         64799    :	result = 16'd12;
         64800    :	result = 16'd12;
         64801    :	result = 16'd13;
         64802    :	result = 16'd13;
         64803    :	result = 16'd13;
         64804    :	result = 16'd13;
         64805    :	result = 16'd13;
         64806    :	result = 16'd13;
         64807    :	result = 16'd13;
         64808    :	result = 16'd13;
         64809    :	result = 16'd13;
         64810    :	result = 16'd13;
         64811    :	result = 16'd13;
         64812    :	result = 16'd13;
         64813    :	result = 16'd13;
         64814    :	result = 16'd13;
         64815    :	result = 16'd13;
         64816    :	result = 16'd13;
         64817    :	result = 16'd13;
         64818    :	result = 16'd13;
         64819    :	result = 16'd13;
         64820    :	result = 16'd13;
         64821    :	result = 16'd13;
         64822    :	result = 16'd14;
         64823    :	result = 16'd14;
         64824    :	result = 16'd14;
         64825    :	result = 16'd14;
         64826    :	result = 16'd14;
         64827    :	result = 16'd14;
         64828    :	result = 16'd14;
         64829    :	result = 16'd14;
         64830    :	result = 16'd14;
         64831    :	result = 16'd14;
         64832    :	result = 16'd14;
         64833    :	result = 16'd14;
         64834    :	result = 16'd14;
         64835    :	result = 16'd14;
         64836    :	result = 16'd14;
         64837    :	result = 16'd14;
         64838    :	result = 16'd14;
         64839    :	result = 16'd14;
         64840    :	result = 16'd14;
         64841    :	result = 16'd14;
         64842    :	result = 16'd15;
         64843    :	result = 16'd15;
         64844    :	result = 16'd15;
         64845    :	result = 16'd15;
         64846    :	result = 16'd15;
         64847    :	result = 16'd15;
         64848    :	result = 16'd15;
         64849    :	result = 16'd15;
         64850    :	result = 16'd15;
         64851    :	result = 16'd15;
         64852    :	result = 16'd15;
         64853    :	result = 16'd15;
         64854    :	result = 16'd15;
         64855    :	result = 16'd15;
         64856    :	result = 16'd15;
         64857    :	result = 16'd15;
         64858    :	result = 16'd15;
         64859    :	result = 16'd15;
         64860    :	result = 16'd15;
         64861    :	result = 16'd16;
         64862    :	result = 16'd16;
         64863    :	result = 16'd16;
         64864    :	result = 16'd16;
         64865    :	result = 16'd16;
         64866    :	result = 16'd16;
         64867    :	result = 16'd16;
         64868    :	result = 16'd16;
         64869    :	result = 16'd16;
         64870    :	result = 16'd16;
         64871    :	result = 16'd16;
         64872    :	result = 16'd16;
         64873    :	result = 16'd16;
         64874    :	result = 16'd16;
         64875    :	result = 16'd16;
         64876    :	result = 16'd16;
         64877    :	result = 16'd16;
         64878    :	result = 16'd16;
         64879    :	result = 16'd17;
         64880    :	result = 16'd17;
         64881    :	result = 16'd17;
         64882    :	result = 16'd17;
         64883    :	result = 16'd17;
         64884    :	result = 16'd17;
         64885    :	result = 16'd17;
         64886    :	result = 16'd17;
         64887    :	result = 16'd17;
         64888    :	result = 16'd17;
         64889    :	result = 16'd17;
         64890    :	result = 16'd17;
         64891    :	result = 16'd17;
         64892    :	result = 16'd17;
         64893    :	result = 16'd17;
         64894    :	result = 16'd17;
         64895    :	result = 16'd17;
         64896    :	result = 16'd18;
         64897    :	result = 16'd18;
         64898    :	result = 16'd18;
         64899    :	result = 16'd18;
         64900    :	result = 16'd18;
         64901    :	result = 16'd18;
         64902    :	result = 16'd18;
         64903    :	result = 16'd18;
         64904    :	result = 16'd18;
         64905    :	result = 16'd18;
         64906    :	result = 16'd18;
         64907    :	result = 16'd18;
         64908    :	result = 16'd18;
         64909    :	result = 16'd18;
         64910    :	result = 16'd18;
         64911    :	result = 16'd18;
         64912    :	result = 16'd18;
         64913    :	result = 16'd19;
         64914    :	result = 16'd19;
         64915    :	result = 16'd19;
         64916    :	result = 16'd19;
         64917    :	result = 16'd19;
         64918    :	result = 16'd19;
         64919    :	result = 16'd19;
         64920    :	result = 16'd19;
         64921    :	result = 16'd19;
         64922    :	result = 16'd19;
         64923    :	result = 16'd19;
         64924    :	result = 16'd19;
         64925    :	result = 16'd19;
         64926    :	result = 16'd19;
         64927    :	result = 16'd19;
         64928    :	result = 16'd19;
         64929    :	result = 16'd20;
         64930    :	result = 16'd20;
         64931    :	result = 16'd20;
         64932    :	result = 16'd20;
         64933    :	result = 16'd20;
         64934    :	result = 16'd20;
         64935    :	result = 16'd20;
         64936    :	result = 16'd20;
         64937    :	result = 16'd20;
         64938    :	result = 16'd20;
         64939    :	result = 16'd20;
         64940    :	result = 16'd20;
         64941    :	result = 16'd20;
         64942    :	result = 16'd20;
         64943    :	result = 16'd20;
         64944    :	result = 16'd21;
         64945    :	result = 16'd21;
         64946    :	result = 16'd21;
         64947    :	result = 16'd21;
         64948    :	result = 16'd21;
         64949    :	result = 16'd21;
         64950    :	result = 16'd21;
         64951    :	result = 16'd21;
         64952    :	result = 16'd21;
         64953    :	result = 16'd21;
         64954    :	result = 16'd21;
         64955    :	result = 16'd21;
         64956    :	result = 16'd21;
         64957    :	result = 16'd21;
         64958    :	result = 16'd22;
         64959    :	result = 16'd22;
         64960    :	result = 16'd22;
         64961    :	result = 16'd22;
         64962    :	result = 16'd22;
         64963    :	result = 16'd22;
         64964    :	result = 16'd22;
         64965    :	result = 16'd22;
         64966    :	result = 16'd22;
         64967    :	result = 16'd22;
         64968    :	result = 16'd22;
         64969    :	result = 16'd22;
         64970    :	result = 16'd22;
         64971    :	result = 16'd22;
         64972    :	result = 16'd23;
         64973    :	result = 16'd23;
         64974    :	result = 16'd23;
         64975    :	result = 16'd23;
         64976    :	result = 16'd23;
         64977    :	result = 16'd23;
         64978    :	result = 16'd23;
         64979    :	result = 16'd23;
         64980    :	result = 16'd23;
         64981    :	result = 16'd23;
         64982    :	result = 16'd23;
         64983    :	result = 16'd23;
         64984    :	result = 16'd23;
         64985    :	result = 16'd23;
         64986    :	result = 16'd24;
         64987    :	result = 16'd24;
         64988    :	result = 16'd24;
         64989    :	result = 16'd24;
         64990    :	result = 16'd24;
         64991    :	result = 16'd24;
         64992    :	result = 16'd24;
         64993    :	result = 16'd24;
         64994    :	result = 16'd24;
         64995    :	result = 16'd24;
         64996    :	result = 16'd24;
         64997    :	result = 16'd24;
         64998    :	result = 16'd24;
         64999    :	result = 16'd25;
         65000    :	result = 16'd25;
         65001    :	result = 16'd25;
         65002    :	result = 16'd25;
         65003    :	result = 16'd25;
         65004    :	result = 16'd25;
         65005    :	result = 16'd25;
         65006    :	result = 16'd25;
         65007    :	result = 16'd25;
         65008    :	result = 16'd25;
         65009    :	result = 16'd25;
         65010    :	result = 16'd25;
         65011    :	result = 16'd25;
         65012    :	result = 16'd26;
         65013    :	result = 16'd26;
         65014    :	result = 16'd26;
         65015    :	result = 16'd26;
         65016    :	result = 16'd26;
         65017    :	result = 16'd26;
         65018    :	result = 16'd26;
         65019    :	result = 16'd26;
         65020    :	result = 16'd26;
         65021    :	result = 16'd26;
         65022    :	result = 16'd26;
         65023    :	result = 16'd26;
         65024    :	result = 16'd26;
         65025    :	result = 16'd27;
         65026    :	result = 16'd27;
         65027    :	result = 16'd27;
         65028    :	result = 16'd27;
         65029    :	result = 16'd27;
         65030    :	result = 16'd27;
         65031    :	result = 16'd27;
         65032    :	result = 16'd27;
         65033    :	result = 16'd27;
         65034    :	result = 16'd27;
         65035    :	result = 16'd27;
         65036    :	result = 16'd27;
         65037    :	result = 16'd28;
         65038    :	result = 16'd28;
         65039    :	result = 16'd28;
         65040    :	result = 16'd28;
         65041    :	result = 16'd28;
         65042    :	result = 16'd28;
         65043    :	result = 16'd28;
         65044    :	result = 16'd28;
         65045    :	result = 16'd28;
         65046    :	result = 16'd28;
         65047    :	result = 16'd28;
         65048    :	result = 16'd28;
         65049    :	result = 16'd29;
         65050    :	result = 16'd29;
         65051    :	result = 16'd29;
         65052    :	result = 16'd29;
         65053    :	result = 16'd29;
         65054    :	result = 16'd29;
         65055    :	result = 16'd29;
         65056    :	result = 16'd29;
         65057    :	result = 16'd29;
         65058    :	result = 16'd29;
         65059    :	result = 16'd29;
         65060    :	result = 16'd29;
         65061    :	result = 16'd30;
         65062    :	result = 16'd30;
         65063    :	result = 16'd30;
         65064    :	result = 16'd30;
         65065    :	result = 16'd30;
         65066    :	result = 16'd30;
         65067    :	result = 16'd30;
         65068    :	result = 16'd30;
         65069    :	result = 16'd30;
         65070    :	result = 16'd30;
         65071    :	result = 16'd30;
         65072    :	result = 16'd30;
         65073    :	result = 16'd31;
         65074    :	result = 16'd31;
         65075    :	result = 16'd31;
         65076    :	result = 16'd31;
         65077    :	result = 16'd31;
         65078    :	result = 16'd31;
         65079    :	result = 16'd31;
         65080    :	result = 16'd31;
         65081    :	result = 16'd31;
         65082    :	result = 16'd31;
         65083    :	result = 16'd31;
         65084    :	result = 16'd32;
         65085    :	result = 16'd32;
         65086    :	result = 16'd32;
         65087    :	result = 16'd32;
         65088    :	result = 16'd32;
         65089    :	result = 16'd32;
         65090    :	result = 16'd32;
         65091    :	result = 16'd32;
         65092    :	result = 16'd32;
         65093    :	result = 16'd32;
         65094    :	result = 16'd32;
         65095    :	result = 16'd33;
         65096    :	result = 16'd33;
         65097    :	result = 16'd33;
         65098    :	result = 16'd33;
         65099    :	result = 16'd33;
         65100    :	result = 16'd33;
         65101    :	result = 16'd33;
         65102    :	result = 16'd33;
         65103    :	result = 16'd33;
         65104    :	result = 16'd33;
         65105    :	result = 16'd33;
         65106    :	result = 16'd33;
         65107    :	result = 16'd34;
         65108    :	result = 16'd34;
         65109    :	result = 16'd34;
         65110    :	result = 16'd34;
         65111    :	result = 16'd34;
         65112    :	result = 16'd34;
         65113    :	result = 16'd34;
         65114    :	result = 16'd34;
         65115    :	result = 16'd34;
         65116    :	result = 16'd34;
         65117    :	result = 16'd35;
         65118    :	result = 16'd35;
         65119    :	result = 16'd35;
         65120    :	result = 16'd35;
         65121    :	result = 16'd35;
         65122    :	result = 16'd35;
         65123    :	result = 16'd35;
         65124    :	result = 16'd35;
         65125    :	result = 16'd35;
         65126    :	result = 16'd35;
         65127    :	result = 16'd35;
         65128    :	result = 16'd36;
         65129    :	result = 16'd36;
         65130    :	result = 16'd36;
         65131    :	result = 16'd36;
         65132    :	result = 16'd36;
         65133    :	result = 16'd36;
         65134    :	result = 16'd36;
         65135    :	result = 16'd36;
         65136    :	result = 16'd36;
         65137    :	result = 16'd36;
         65138    :	result = 16'd36;
         65139    :	result = 16'd37;
         65140    :	result = 16'd37;
         65141    :	result = 16'd37;
         65142    :	result = 16'd37;
         65143    :	result = 16'd37;
         65144    :	result = 16'd37;
         65145    :	result = 16'd37;
         65146    :	result = 16'd37;
         65147    :	result = 16'd37;
         65148    :	result = 16'd37;
         65149    :	result = 16'd37;
         65150    :	result = 16'd38;
         65151    :	result = 16'd38;
         65152    :	result = 16'd38;
         65153    :	result = 16'd38;
         65154    :	result = 16'd38;
         65155    :	result = 16'd38;
         65156    :	result = 16'd38;
         65157    :	result = 16'd38;
         65158    :	result = 16'd38;
         65159    :	result = 16'd38;
         65160    :	result = 16'd39;
         65161    :	result = 16'd39;
         65162    :	result = 16'd39;
         65163    :	result = 16'd39;
         65164    :	result = 16'd39;
         65165    :	result = 16'd39;
         65166    :	result = 16'd39;
         65167    :	result = 16'd39;
         65168    :	result = 16'd39;
         65169    :	result = 16'd39;
         65170    :	result = 16'd39;
         65171    :	result = 16'd40;
         65172    :	result = 16'd40;
         65173    :	result = 16'd40;
         65174    :	result = 16'd40;
         65175    :	result = 16'd40;
         65176    :	result = 16'd40;
         65177    :	result = 16'd40;
         65178    :	result = 16'd40;
         65179    :	result = 16'd40;
         65180    :	result = 16'd40;
         65181    :	result = 16'd41;
         65182    :	result = 16'd41;
         65183    :	result = 16'd41;
         65184    :	result = 16'd41;
         65185    :	result = 16'd41;
         65186    :	result = 16'd41;
         65187    :	result = 16'd41;
         65188    :	result = 16'd41;
         65189    :	result = 16'd41;
         65190    :	result = 16'd41;
         65191    :	result = 16'd42;
         65192    :	result = 16'd42;
         65193    :	result = 16'd42;
         65194    :	result = 16'd42;
         65195    :	result = 16'd42;
         65196    :	result = 16'd42;
         65197    :	result = 16'd42;
         65198    :	result = 16'd42;
         65199    :	result = 16'd42;
         65200    :	result = 16'd42;
         65201    :	result = 16'd42;
         65202    :	result = 16'd43;
         65203    :	result = 16'd43;
         65204    :	result = 16'd43;
         65205    :	result = 16'd43;
         65206    :	result = 16'd43;
         65207    :	result = 16'd43;
         65208    :	result = 16'd43;
         65209    :	result = 16'd43;
         65210    :	result = 16'd43;
         65211    :	result = 16'd43;
         65212    :	result = 16'd44;
         65213    :	result = 16'd44;
         65214    :	result = 16'd44;
         65215    :	result = 16'd44;
         65216    :	result = 16'd44;
         65217    :	result = 16'd44;
         65218    :	result = 16'd44;
         65219    :	result = 16'd44;
         65220    :	result = 16'd44;
         65221    :	result = 16'd44;
         65222    :	result = 16'd44;
         65223    :	result = 16'd45;
         65224    :	result = 16'd45;
         65225    :	result = 16'd45;
         65226    :	result = 16'd45;
         65227    :	result = 16'd45;
         65228    :	result = 16'd45;
         65229    :	result = 16'd45;
         65230    :	result = 16'd45;
         65231    :	result = 16'd45;
         65232    :	result = 16'd45;
         65233    :	result = 16'd46;
         65234    :	result = 16'd46;
         65235    :	result = 16'd46;
         65236    :	result = 16'd46;
         65237    :	result = 16'd46;
         65238    :	result = 16'd46;
         65239    :	result = 16'd46;
         65240    :	result = 16'd46;
         65241    :	result = 16'd46;
         65242    :	result = 16'd46;
         65243    :	result = 16'd46;
         65244    :	result = 16'd47;
         65245    :	result = 16'd47;
         65246    :	result = 16'd47;
         65247    :	result = 16'd47;
         65248    :	result = 16'd47;
         65249    :	result = 16'd47;
         65250    :	result = 16'd47;
         65251    :	result = 16'd47;
         65252    :	result = 16'd47;
         65253    :	result = 16'd47;
         65254    :	result = 16'd48;
         65255    :	result = 16'd48;
         65256    :	result = 16'd48;
         65257    :	result = 16'd48;
         65258    :	result = 16'd48;
         65259    :	result = 16'd48;
         65260    :	result = 16'd48;
         65261    :	result = 16'd48;
         65262    :	result = 16'd48;
         65263    :	result = 16'd48;
         65264    :	result = 16'd48;
         65265    :	result = 16'd49;
         65266    :	result = 16'd49;
         65267    :	result = 16'd49;
         65268    :	result = 16'd49;
         65269    :	result = 16'd49;
         65270    :	result = 16'd49;
         65271    :	result = 16'd49;
         65272    :	result = 16'd49;
         65273    :	result = 16'd49;
         65274    :	result = 16'd49;
         65275    :	result = 16'd49;
         65276    :	result = 16'd50;
         65277    :	result = 16'd50;
         65278    :	result = 16'd50;
         65279    :	result = 16'd50;
         65280    :	result = 16'd50;
         65281    :	result = 16'd50;
         65282    :	result = 16'd50;
         65283    :	result = 16'd50;
         65284    :	result = 16'd50;
         65285    :	result = 16'd50;
         65286    :	result = 16'd50;
         65287    :	result = 16'd51;
         65288    :	result = 16'd51;
         65289    :	result = 16'd51;
         65290    :	result = 16'd51;
         65291    :	result = 16'd51;
         65292    :	result = 16'd51;
         65293    :	result = 16'd51;
         65294    :	result = 16'd51;
         65295    :	result = 16'd51;
         65296    :	result = 16'd51;
         65297    :	result = 16'd51;
         65298    :	result = 16'd52;
         65299    :	result = 16'd52;
         65300    :	result = 16'd52;
         65301    :	result = 16'd52;
         65302    :	result = 16'd52;
         65303    :	result = 16'd52;
         65304    :	result = 16'd52;
         65305    :	result = 16'd52;
         65306    :	result = 16'd52;
         65307    :	result = 16'd52;
         65308    :	result = 16'd52;
         65309    :	result = 16'd52;
         65310    :	result = 16'd53;
         65311    :	result = 16'd53;
         65312    :	result = 16'd53;
         65313    :	result = 16'd53;
         65314    :	result = 16'd53;
         65315    :	result = 16'd53;
         65316    :	result = 16'd53;
         65317    :	result = 16'd53;
         65318    :	result = 16'd53;
         65319    :	result = 16'd53;
         65320    :	result = 16'd53;
         65321    :	result = 16'd54;
         65322    :	result = 16'd54;
         65323    :	result = 16'd54;
         65324    :	result = 16'd54;
         65325    :	result = 16'd54;
         65326    :	result = 16'd54;
         65327    :	result = 16'd54;
         65328    :	result = 16'd54;
         65329    :	result = 16'd54;
         65330    :	result = 16'd54;
         65331    :	result = 16'd54;
         65332    :	result = 16'd54;
         65333    :	result = 16'd54;
         65334    :	result = 16'd55;
         65335    :	result = 16'd55;
         65336    :	result = 16'd55;
         65337    :	result = 16'd55;
         65338    :	result = 16'd55;
         65339    :	result = 16'd55;
         65340    :	result = 16'd55;
         65341    :	result = 16'd55;
         65342    :	result = 16'd55;
         65343    :	result = 16'd55;
         65344    :	result = 16'd55;
         65345    :	result = 16'd55;
         65346    :	result = 16'd56;
         65347    :	result = 16'd56;
         65348    :	result = 16'd56;
         65349    :	result = 16'd56;
         65350    :	result = 16'd56;
         65351    :	result = 16'd56;
         65352    :	result = 16'd56;
         65353    :	result = 16'd56;
         65354    :	result = 16'd56;
         65355    :	result = 16'd56;
         65356    :	result = 16'd56;
         65357    :	result = 16'd56;
         65358    :	result = 16'd56;
         65359    :	result = 16'd56;
         65360    :	result = 16'd57;
         65361    :	result = 16'd57;
         65362    :	result = 16'd57;
         65363    :	result = 16'd57;
         65364    :	result = 16'd57;
         65365    :	result = 16'd57;
         65366    :	result = 16'd57;
         65367    :	result = 16'd57;
         65368    :	result = 16'd57;
         65369    :	result = 16'd57;
         65370    :	result = 16'd57;
         65371    :	result = 16'd57;
         65372    :	result = 16'd57;
         65373    :	result = 16'd57;
         65374    :	result = 16'd58;
         65375    :	result = 16'd58;
         65376    :	result = 16'd58;
         65377    :	result = 16'd58;
         65378    :	result = 16'd58;
         65379    :	result = 16'd58;
         65380    :	result = 16'd58;
         65381    :	result = 16'd58;
         65382    :	result = 16'd58;
         65383    :	result = 16'd58;
         65384    :	result = 16'd58;
         65385    :	result = 16'd58;
         65386    :	result = 16'd58;
         65387    :	result = 16'd58;
         65388    :	result = 16'd59;
         65389    :	result = 16'd59;
         65390    :	result = 16'd59;
         65391    :	result = 16'd59;
         65392    :	result = 16'd59;
         65393    :	result = 16'd59;
         65394    :	result = 16'd59;
         65395    :	result = 16'd59;
         65396    :	result = 16'd59;
         65397    :	result = 16'd59;
         65398    :	result = 16'd59;
         65399    :	result = 16'd59;
         65400    :	result = 16'd59;
         65401    :	result = 16'd59;
         65402    :	result = 16'd59;
         65403    :	result = 16'd59;
         65404    :	result = 16'd59;
         65405    :	result = 16'd60;
         65406    :	result = 16'd60;
         65407    :	result = 16'd60;
         65408    :	result = 16'd60;
         65409    :	result = 16'd60;
         65410    :	result = 16'd60;
         65411    :	result = 16'd60;
         65412    :	result = 16'd60;
         65413    :	result = 16'd60;
         65414    :	result = 16'd60;
         65415    :	result = 16'd60;
         65416    :	result = 16'd60;
         65417    :	result = 16'd60;
         65418    :	result = 16'd60;
         65419    :	result = 16'd60;
         65420    :	result = 16'd60;
         65421    :	result = 16'd60;
         65422    :	result = 16'd60;
         65423    :	result = 16'd61;
         65424    :	result = 16'd61;
         65425    :	result = 16'd61;
         65426    :	result = 16'd61;
         65427    :	result = 16'd61;
         65428    :	result = 16'd61;
         65429    :	result = 16'd61;
         65430    :	result = 16'd61;
         65431    :	result = 16'd61;
         65432    :	result = 16'd61;
         65433    :	result = 16'd61;
         65434    :	result = 16'd61;
         65435    :	result = 16'd61;
         65436    :	result = 16'd61;
         65437    :	result = 16'd61;
         65438    :	result = 16'd61;
         65439    :	result = 16'd61;
         65440    :	result = 16'd61;
         65441    :	result = 16'd61;
         65442    :	result = 16'd61;
         65443    :	result = 16'd61;
         65444    :	result = 16'd62;
         65445    :	result = 16'd62;
         65446    :	result = 16'd62;
         65447    :	result = 16'd62;
         65448    :	result = 16'd62;
         65449    :	result = 16'd62;
         65450    :	result = 16'd62;
         65451    :	result = 16'd62;
         65452    :	result = 16'd62;
         65453    :	result = 16'd62;
         65454    :	result = 16'd62;
         65455    :	result = 16'd62;
         65456    :	result = 16'd62;
         65457    :	result = 16'd62;
         65458    :	result = 16'd62;
         65459    :	result = 16'd62;
         65460    :	result = 16'd62;
         65461    :	result = 16'd62;
         65462    :	result = 16'd62;
         65463    :	result = 16'd62;
         65464    :	result = 16'd62;
         65465    :	result = 16'd62;
         65466    :	result = 16'd62;
         65467    :	result = 16'd62;
         65468    :	result = 16'd62;
         65469    :	result = 16'd62;
         65470    :	result = 16'd62;
         65471    :	result = 16'd63;
         65472    :	result = 16'd63;
         65473    :	result = 16'd63;
         65474    :	result = 16'd63;
         65475    :	result = 16'd63;
         65476    :	result = 16'd63;
         65477    :	result = 16'd63;
         65478    :	result = 16'd63;
         65479    :	result = 16'd63;
         65480    :	result = 16'd63;
         65481    :	result = 16'd63;
         65482    :	result = 16'd63;
         65483    :	result = 16'd63;
         65484    :	result = 16'd63;
         65485    :	result = 16'd63;
         65486    :	result = 16'd63;
         65487    :	result = 16'd63;
         65488    :	result = 16'd63;
         65489    :	result = 16'd63;
         65490    :	result = 16'd63;
         65491    :	result = 16'd63;
         65492    :	result = 16'd63;
         65493    :	result = 16'd63;
         65494    :	result = 16'd63;
         65495    :	result = 16'd63;
         65496    :	result = 16'd63;
         65497    :	result = 16'd63;
         65498    :	result = 16'd63;
         65499    :	result = 16'd63;
         65500    :	result = 16'd63;
         65501    :	result = 16'd63;
         65502    :	result = 16'd63;
         65503    :	result = 16'd63;
         65504    :	result = 16'd63;
         65505    :	result = 16'd63;
         65506    :	result = 16'd63;
         65507    :	result = 16'd63;
         65508    :	result = 16'd63;
         65509    :	result = 16'd63;
         65510    :	result = 16'd63;
         65511    :	result = 16'd63;
         65512    :	result = 16'd63;
         65513    :	result = 16'd63;
         65514    :	result = 16'd63;
         65515    :	result = 16'd63;
         65516    :	result = 16'd63;
         65517    :	result = 16'd63;
         65518    :	result = 16'd63;
         65519    :	result = 16'd63;
         65520    :	result = 16'd63;
         65521    :	result = 16'd63;
         65522    :	result = 16'd63;
         65523    :	result = 16'd63;
         65524    :	result = 16'd63;
         65525    :	result = 16'd63;
         65526    :	result = 16'd63;
         65527    :	result = 16'd63;
         65528    :	result = 16'd63;
         65529    :	result = 16'd63;
         65530    :	result = 16'd63;
         65531    :	result = 16'd63;
         65532    :	result = 16'd63;
         65533    :	result = 16'd63;
         65534    :	result = 16'd63;
         65535    :	result = 16'd64;
         0        :	result = 16'd63;
         1        :	result = 16'd63;
         2        :	result = 16'd63;
         3        :	result = 16'd63;
         4        :	result = 16'd63;
         5        :	result = 16'd63;
         6        :	result = 16'd63;
         7        :	result = 16'd63;
         8        :	result = 16'd63;
         9        :	result = 16'd63;
         10       :	result = 16'd63;
         11       :	result = 16'd63;
         12       :	result = 16'd63;
         13       :	result = 16'd63;
         14       :	result = 16'd63;
         15       :	result = 16'd63;
         16       :	result = 16'd63;
         17       :	result = 16'd63;
         18       :	result = 16'd63;
         19       :	result = 16'd63;
         20       :	result = 16'd63;
         21       :	result = 16'd63;
         22       :	result = 16'd63;
         23       :	result = 16'd63;
         24       :	result = 16'd63;
         25       :	result = 16'd63;
         26       :	result = 16'd63;
         27       :	result = 16'd63;
         28       :	result = 16'd63;
         29       :	result = 16'd63;
         30       :	result = 16'd63;
         31       :	result = 16'd63;
         32       :	result = 16'd63;
         33       :	result = 16'd63;
         34       :	result = 16'd63;
         35       :	result = 16'd63;
         36       :	result = 16'd63;
         37       :	result = 16'd63;
         38       :	result = 16'd63;
         39       :	result = 16'd63;
         40       :	result = 16'd63;
         41       :	result = 16'd63;
         42       :	result = 16'd63;
         43       :	result = 16'd63;
         44       :	result = 16'd63;
         45       :	result = 16'd63;
         46       :	result = 16'd63;
         47       :	result = 16'd63;
         48       :	result = 16'd63;
         49       :	result = 16'd63;
         50       :	result = 16'd63;
         51       :	result = 16'd63;
         52       :	result = 16'd63;
         53       :	result = 16'd63;
         54       :	result = 16'd63;
         55       :	result = 16'd63;
         56       :	result = 16'd63;
         57       :	result = 16'd63;
         58       :	result = 16'd63;
         59       :	result = 16'd63;
         60       :	result = 16'd63;
         61       :	result = 16'd63;
         62       :	result = 16'd63;
         63       :	result = 16'd63;
         64       :	result = 16'd62;
         65       :	result = 16'd62;
         66       :	result = 16'd62;
         67       :	result = 16'd62;
         68       :	result = 16'd62;
         69       :	result = 16'd62;
         70       :	result = 16'd62;
         71       :	result = 16'd62;
         72       :	result = 16'd62;
         73       :	result = 16'd62;
         74       :	result = 16'd62;
         75       :	result = 16'd62;
         76       :	result = 16'd62;
         77       :	result = 16'd62;
         78       :	result = 16'd62;
         79       :	result = 16'd62;
         80       :	result = 16'd62;
         81       :	result = 16'd62;
         82       :	result = 16'd62;
         83       :	result = 16'd62;
         84       :	result = 16'd62;
         85       :	result = 16'd62;
         86       :	result = 16'd62;
         87       :	result = 16'd62;
         88       :	result = 16'd62;
         89       :	result = 16'd62;
         90       :	result = 16'd62;
         91       :	result = 16'd61;
         92       :	result = 16'd61;
         93       :	result = 16'd61;
         94       :	result = 16'd61;
         95       :	result = 16'd61;
         96       :	result = 16'd61;
         97       :	result = 16'd61;
         98       :	result = 16'd61;
         99       :	result = 16'd61;
         100      :	result = 16'd61;
         101      :	result = 16'd61;
         102      :	result = 16'd61;
         103      :	result = 16'd61;
         104      :	result = 16'd61;
         105      :	result = 16'd61;
         106      :	result = 16'd61;
         107      :	result = 16'd61;
         108      :	result = 16'd61;
         109      :	result = 16'd61;
         110      :	result = 16'd61;
         111      :	result = 16'd61;
         112      :	result = 16'd60;
         113      :	result = 16'd60;
         114      :	result = 16'd60;
         115      :	result = 16'd60;
         116      :	result = 16'd60;
         117      :	result = 16'd60;
         118      :	result = 16'd60;
         119      :	result = 16'd60;
         120      :	result = 16'd60;
         121      :	result = 16'd60;
         122      :	result = 16'd60;
         123      :	result = 16'd60;
         124      :	result = 16'd60;
         125      :	result = 16'd60;
         126      :	result = 16'd60;
         127      :	result = 16'd60;
         128      :	result = 16'd60;
         129      :	result = 16'd60;
         130      :	result = 16'd59;
         131      :	result = 16'd59;
         132      :	result = 16'd59;
         133      :	result = 16'd59;
         134      :	result = 16'd59;
         135      :	result = 16'd59;
         136      :	result = 16'd59;
         137      :	result = 16'd59;
         138      :	result = 16'd59;
         139      :	result = 16'd59;
         140      :	result = 16'd59;
         141      :	result = 16'd59;
         142      :	result = 16'd59;
         143      :	result = 16'd59;
         144      :	result = 16'd59;
         145      :	result = 16'd59;
         146      :	result = 16'd59;
         147      :	result = 16'd58;
         148      :	result = 16'd58;
         149      :	result = 16'd58;
         150      :	result = 16'd58;
         151      :	result = 16'd58;
         152      :	result = 16'd58;
         153      :	result = 16'd58;
         154      :	result = 16'd58;
         155      :	result = 16'd58;
         156      :	result = 16'd58;
         157      :	result = 16'd58;
         158      :	result = 16'd58;
         159      :	result = 16'd58;
         160      :	result = 16'd58;
         161      :	result = 16'd57;
         162      :	result = 16'd57;
         163      :	result = 16'd57;
         164      :	result = 16'd57;
         165      :	result = 16'd57;
         166      :	result = 16'd57;
         167      :	result = 16'd57;
         168      :	result = 16'd57;
         169      :	result = 16'd57;
         170      :	result = 16'd57;
         171      :	result = 16'd57;
         172      :	result = 16'd57;
         173      :	result = 16'd57;
         174      :	result = 16'd57;
         175      :	result = 16'd56;
         176      :	result = 16'd56;
         177      :	result = 16'd56;
         178      :	result = 16'd56;
         179      :	result = 16'd56;
         180      :	result = 16'd56;
         181      :	result = 16'd56;
         182      :	result = 16'd56;
         183      :	result = 16'd56;
         184      :	result = 16'd56;
         185      :	result = 16'd56;
         186      :	result = 16'd56;
         187      :	result = 16'd56;
         188      :	result = 16'd56;
         189      :	result = 16'd55;
         190      :	result = 16'd55;
         191      :	result = 16'd55;
         192      :	result = 16'd55;
         193      :	result = 16'd55;
         194      :	result = 16'd55;
         195      :	result = 16'd55;
         196      :	result = 16'd55;
         197      :	result = 16'd55;
         198      :	result = 16'd55;
         199      :	result = 16'd55;
         200      :	result = 16'd55;
         201      :	result = 16'd54;
         202      :	result = 16'd54;
         203      :	result = 16'd54;
         204      :	result = 16'd54;
         205      :	result = 16'd54;
         206      :	result = 16'd54;
         207      :	result = 16'd54;
         208      :	result = 16'd54;
         209      :	result = 16'd54;
         210      :	result = 16'd54;
         211      :	result = 16'd54;
         212      :	result = 16'd54;
         213      :	result = 16'd54;
         214      :	result = 16'd53;
         215      :	result = 16'd53;
         216      :	result = 16'd53;
         217      :	result = 16'd53;
         218      :	result = 16'd53;
         219      :	result = 16'd53;
         220      :	result = 16'd53;
         221      :	result = 16'd53;
         222      :	result = 16'd53;
         223      :	result = 16'd53;
         224      :	result = 16'd53;
         225      :	result = 16'd52;
         226      :	result = 16'd52;
         227      :	result = 16'd52;
         228      :	result = 16'd52;
         229      :	result = 16'd52;
         230      :	result = 16'd52;
         231      :	result = 16'd52;
         232      :	result = 16'd52;
         233      :	result = 16'd52;
         234      :	result = 16'd52;
         235      :	result = 16'd52;
         236      :	result = 16'd52;
         237      :	result = 16'd51;
         238      :	result = 16'd51;
         239      :	result = 16'd51;
         240      :	result = 16'd51;
         241      :	result = 16'd51;
         242      :	result = 16'd51;
         243      :	result = 16'd51;
         244      :	result = 16'd51;
         245      :	result = 16'd51;
         246      :	result = 16'd51;
         247      :	result = 16'd51;
         248      :	result = 16'd50;
         249      :	result = 16'd50;
         250      :	result = 16'd50;
         251      :	result = 16'd50;
         252      :	result = 16'd50;
         253      :	result = 16'd50;
         254      :	result = 16'd50;
         255      :	result = 16'd50;
         256      :	result = 16'd50;
         257      :	result = 16'd50;
         258      :	result = 16'd50;
         259      :	result = 16'd49;
         260      :	result = 16'd49;
         261      :	result = 16'd49;
         262      :	result = 16'd49;
         263      :	result = 16'd49;
         264      :	result = 16'd49;
         265      :	result = 16'd49;
         266      :	result = 16'd49;
         267      :	result = 16'd49;
         268      :	result = 16'd49;
         269      :	result = 16'd49;
         270      :	result = 16'd48;
         271      :	result = 16'd48;
         272      :	result = 16'd48;
         273      :	result = 16'd48;
         274      :	result = 16'd48;
         275      :	result = 16'd48;
         276      :	result = 16'd48;
         277      :	result = 16'd48;
         278      :	result = 16'd48;
         279      :	result = 16'd48;
         280      :	result = 16'd48;
         281      :	result = 16'd47;
         282      :	result = 16'd47;
         283      :	result = 16'd47;
         284      :	result = 16'd47;
         285      :	result = 16'd47;
         286      :	result = 16'd47;
         287      :	result = 16'd47;
         288      :	result = 16'd47;
         289      :	result = 16'd47;
         290      :	result = 16'd47;
         291      :	result = 16'd46;
         292      :	result = 16'd46;
         293      :	result = 16'd46;
         294      :	result = 16'd46;
         295      :	result = 16'd46;
         296      :	result = 16'd46;
         297      :	result = 16'd46;
         298      :	result = 16'd46;
         299      :	result = 16'd46;
         300      :	result = 16'd46;
         301      :	result = 16'd46;
         302      :	result = 16'd45;
         303      :	result = 16'd45;
         304      :	result = 16'd45;
         305      :	result = 16'd45;
         306      :	result = 16'd45;
         307      :	result = 16'd45;
         308      :	result = 16'd45;
         309      :	result = 16'd45;
         310      :	result = 16'd45;
         311      :	result = 16'd45;
         312      :	result = 16'd44;
         313      :	result = 16'd44;
         314      :	result = 16'd44;
         315      :	result = 16'd44;
         316      :	result = 16'd44;
         317      :	result = 16'd44;
         318      :	result = 16'd44;
         319      :	result = 16'd44;
         320      :	result = 16'd44;
         321      :	result = 16'd44;
         322      :	result = 16'd44;
         323      :	result = 16'd43;
         324      :	result = 16'd43;
         325      :	result = 16'd43;
         326      :	result = 16'd43;
         327      :	result = 16'd43;
         328      :	result = 16'd43;
         329      :	result = 16'd43;
         330      :	result = 16'd43;
         331      :	result = 16'd43;
         332      :	result = 16'd43;
         333      :	result = 16'd42;
         334      :	result = 16'd42;
         335      :	result = 16'd42;
         336      :	result = 16'd42;
         337      :	result = 16'd42;
         338      :	result = 16'd42;
         339      :	result = 16'd42;
         340      :	result = 16'd42;
         341      :	result = 16'd42;
         342      :	result = 16'd42;
         343      :	result = 16'd42;
         344      :	result = 16'd41;
         345      :	result = 16'd41;
         346      :	result = 16'd41;
         347      :	result = 16'd41;
         348      :	result = 16'd41;
         349      :	result = 16'd41;
         350      :	result = 16'd41;
         351      :	result = 16'd41;
         352      :	result = 16'd41;
         353      :	result = 16'd41;
         354      :	result = 16'd40;
         355      :	result = 16'd40;
         356      :	result = 16'd40;
         357      :	result = 16'd40;
         358      :	result = 16'd40;
         359      :	result = 16'd40;
         360      :	result = 16'd40;
         361      :	result = 16'd40;
         362      :	result = 16'd40;
         363      :	result = 16'd40;
         364      :	result = 16'd39;
         365      :	result = 16'd39;
         366      :	result = 16'd39;
         367      :	result = 16'd39;
         368      :	result = 16'd39;
         369      :	result = 16'd39;
         370      :	result = 16'd39;
         371      :	result = 16'd39;
         372      :	result = 16'd39;
         373      :	result = 16'd39;
         374      :	result = 16'd39;
         375      :	result = 16'd38;
         376      :	result = 16'd38;
         377      :	result = 16'd38;
         378      :	result = 16'd38;
         379      :	result = 16'd38;
         380      :	result = 16'd38;
         381      :	result = 16'd38;
         382      :	result = 16'd38;
         383      :	result = 16'd38;
         384      :	result = 16'd38;
         385      :	result = 16'd37;
         386      :	result = 16'd37;
         387      :	result = 16'd37;
         388      :	result = 16'd37;
         389      :	result = 16'd37;
         390      :	result = 16'd37;
         391      :	result = 16'd37;
         392      :	result = 16'd37;
         393      :	result = 16'd37;
         394      :	result = 16'd37;
         395      :	result = 16'd37;
         396      :	result = 16'd36;
         397      :	result = 16'd36;
         398      :	result = 16'd36;
         399      :	result = 16'd36;
         400      :	result = 16'd36;
         401      :	result = 16'd36;
         402      :	result = 16'd36;
         403      :	result = 16'd36;
         404      :	result = 16'd36;
         405      :	result = 16'd36;
         406      :	result = 16'd36;
         407      :	result = 16'd35;
         408      :	result = 16'd35;
         409      :	result = 16'd35;
         410      :	result = 16'd35;
         411      :	result = 16'd35;
         412      :	result = 16'd35;
         413      :	result = 16'd35;
         414      :	result = 16'd35;
         415      :	result = 16'd35;
         416      :	result = 16'd35;
         417      :	result = 16'd35;
         418      :	result = 16'd34;
         419      :	result = 16'd34;
         420      :	result = 16'd34;
         421      :	result = 16'd34;
         422      :	result = 16'd34;
         423      :	result = 16'd34;
         424      :	result = 16'd34;
         425      :	result = 16'd34;
         426      :	result = 16'd34;
         427      :	result = 16'd34;
         428      :	result = 16'd33;
         429      :	result = 16'd33;
         430      :	result = 16'd33;
         431      :	result = 16'd33;
         432      :	result = 16'd33;
         433      :	result = 16'd33;
         434      :	result = 16'd33;
         435      :	result = 16'd33;
         436      :	result = 16'd33;
         437      :	result = 16'd33;
         438      :	result = 16'd33;
         439      :	result = 16'd33;
         440      :	result = 16'd32;
         441      :	result = 16'd32;
         442      :	result = 16'd32;
         443      :	result = 16'd32;
         444      :	result = 16'd32;
         445      :	result = 16'd32;
         446      :	result = 16'd32;
         447      :	result = 16'd32;
         448      :	result = 16'd32;
         449      :	result = 16'd32;
         450      :	result = 16'd32;
         451      :	result = 16'd31;
         452      :	result = 16'd31;
         453      :	result = 16'd31;
         454      :	result = 16'd31;
         455      :	result = 16'd31;
         456      :	result = 16'd31;
         457      :	result = 16'd31;
         458      :	result = 16'd31;
         459      :	result = 16'd31;
         460      :	result = 16'd31;
         461      :	result = 16'd31;
         462      :	result = 16'd30;
         463      :	result = 16'd30;
         464      :	result = 16'd30;
         465      :	result = 16'd30;
         466      :	result = 16'd30;
         467      :	result = 16'd30;
         468      :	result = 16'd30;
         469      :	result = 16'd30;
         470      :	result = 16'd30;
         471      :	result = 16'd30;
         472      :	result = 16'd30;
         473      :	result = 16'd30;
         474      :	result = 16'd29;
         475      :	result = 16'd29;
         476      :	result = 16'd29;
         477      :	result = 16'd29;
         478      :	result = 16'd29;
         479      :	result = 16'd29;
         480      :	result = 16'd29;
         481      :	result = 16'd29;
         482      :	result = 16'd29;
         483      :	result = 16'd29;
         484      :	result = 16'd29;
         485      :	result = 16'd29;
         486      :	result = 16'd28;
         487      :	result = 16'd28;
         488      :	result = 16'd28;
         489      :	result = 16'd28;
         490      :	result = 16'd28;
         491      :	result = 16'd28;
         492      :	result = 16'd28;
         493      :	result = 16'd28;
         494      :	result = 16'd28;
         495      :	result = 16'd28;
         496      :	result = 16'd28;
         497      :	result = 16'd28;
         498      :	result = 16'd27;
         499      :	result = 16'd27;
         500      :	result = 16'd27;
         501      :	result = 16'd27;
         502      :	result = 16'd27;
         503      :	result = 16'd27;
         504      :	result = 16'd27;
         505      :	result = 16'd27;
         506      :	result = 16'd27;
         507      :	result = 16'd27;
         508      :	result = 16'd27;
         509      :	result = 16'd27;
         510      :	result = 16'd26;
         511      :	result = 16'd26;
         512      :	result = 16'd26;
         513      :	result = 16'd26;
         514      :	result = 16'd26;
         515      :	result = 16'd26;
         516      :	result = 16'd26;
         517      :	result = 16'd26;
         518      :	result = 16'd26;
         519      :	result = 16'd26;
         520      :	result = 16'd26;
         521      :	result = 16'd26;
         522      :	result = 16'd26;
         523      :	result = 16'd25;
         524      :	result = 16'd25;
         525      :	result = 16'd25;
         526      :	result = 16'd25;
         527      :	result = 16'd25;
         528      :	result = 16'd25;
         529      :	result = 16'd25;
         530      :	result = 16'd25;
         531      :	result = 16'd25;
         532      :	result = 16'd25;
         533      :	result = 16'd25;
         534      :	result = 16'd25;
         535      :	result = 16'd25;
         536      :	result = 16'd24;
         537      :	result = 16'd24;
         538      :	result = 16'd24;
         539      :	result = 16'd24;
         540      :	result = 16'd24;
         541      :	result = 16'd24;
         542      :	result = 16'd24;
         543      :	result = 16'd24;
         544      :	result = 16'd24;
         545      :	result = 16'd24;
         546      :	result = 16'd24;
         547      :	result = 16'd24;
         548      :	result = 16'd24;
         549      :	result = 16'd23;
         550      :	result = 16'd23;
         551      :	result = 16'd23;
         552      :	result = 16'd23;
         553      :	result = 16'd23;
         554      :	result = 16'd23;
         555      :	result = 16'd23;
         556      :	result = 16'd23;
         557      :	result = 16'd23;
         558      :	result = 16'd23;
         559      :	result = 16'd23;
         560      :	result = 16'd23;
         561      :	result = 16'd23;
         562      :	result = 16'd23;
         563      :	result = 16'd22;
         564      :	result = 16'd22;
         565      :	result = 16'd22;
         566      :	result = 16'd22;
         567      :	result = 16'd22;
         568      :	result = 16'd22;
         569      :	result = 16'd22;
         570      :	result = 16'd22;
         571      :	result = 16'd22;
         572      :	result = 16'd22;
         573      :	result = 16'd22;
         574      :	result = 16'd22;
         575      :	result = 16'd22;
         576      :	result = 16'd22;
         577      :	result = 16'd21;
         578      :	result = 16'd21;
         579      :	result = 16'd21;
         580      :	result = 16'd21;
         581      :	result = 16'd21;
         582      :	result = 16'd21;
         583      :	result = 16'd21;
         584      :	result = 16'd21;
         585      :	result = 16'd21;
         586      :	result = 16'd21;
         587      :	result = 16'd21;
         588      :	result = 16'd21;
         589      :	result = 16'd21;
         590      :	result = 16'd21;
         591      :	result = 16'd20;
         592      :	result = 16'd20;
         593      :	result = 16'd20;
         594      :	result = 16'd20;
         595      :	result = 16'd20;
         596      :	result = 16'd20;
         597      :	result = 16'd20;
         598      :	result = 16'd20;
         599      :	result = 16'd20;
         600      :	result = 16'd20;
         601      :	result = 16'd20;
         602      :	result = 16'd20;
         603      :	result = 16'd20;
         604      :	result = 16'd20;
         605      :	result = 16'd20;
         606      :	result = 16'd19;
         607      :	result = 16'd19;
         608      :	result = 16'd19;
         609      :	result = 16'd19;
         610      :	result = 16'd19;
         611      :	result = 16'd19;
         612      :	result = 16'd19;
         613      :	result = 16'd19;
         614      :	result = 16'd19;
         615      :	result = 16'd19;
         616      :	result = 16'd19;
         617      :	result = 16'd19;
         618      :	result = 16'd19;
         619      :	result = 16'd19;
         620      :	result = 16'd19;
         621      :	result = 16'd19;
         622      :	result = 16'd18;
         623      :	result = 16'd18;
         624      :	result = 16'd18;
         625      :	result = 16'd18;
         626      :	result = 16'd18;
         627      :	result = 16'd18;
         628      :	result = 16'd18;
         629      :	result = 16'd18;
         630      :	result = 16'd18;
         631      :	result = 16'd18;
         632      :	result = 16'd18;
         633      :	result = 16'd18;
         634      :	result = 16'd18;
         635      :	result = 16'd18;
         636      :	result = 16'd18;
         637      :	result = 16'd18;
         638      :	result = 16'd18;
         639      :	result = 16'd17;
         640      :	result = 16'd17;
         641      :	result = 16'd17;
         642      :	result = 16'd17;
         643      :	result = 16'd17;
         644      :	result = 16'd17;
         645      :	result = 16'd17;
         646      :	result = 16'd17;
         647      :	result = 16'd17;
         648      :	result = 16'd17;
         649      :	result = 16'd17;
         650      :	result = 16'd17;
         651      :	result = 16'd17;
         652      :	result = 16'd17;
         653      :	result = 16'd17;
         654      :	result = 16'd17;
         655      :	result = 16'd17;
         656      :	result = 16'd16;
         657      :	result = 16'd16;
         658      :	result = 16'd16;
         659      :	result = 16'd16;
         660      :	result = 16'd16;
         661      :	result = 16'd16;
         662      :	result = 16'd16;
         663      :	result = 16'd16;
         664      :	result = 16'd16;
         665      :	result = 16'd16;
         666      :	result = 16'd16;
         667      :	result = 16'd16;
         668      :	result = 16'd16;
         669      :	result = 16'd16;
         670      :	result = 16'd16;
         671      :	result = 16'd16;
         672      :	result = 16'd16;
         673      :	result = 16'd16;
         674      :	result = 16'd15;
         675      :	result = 16'd15;
         676      :	result = 16'd15;
         677      :	result = 16'd15;
         678      :	result = 16'd15;
         679      :	result = 16'd15;
         680      :	result = 16'd15;
         681      :	result = 16'd15;
         682      :	result = 16'd15;
         683      :	result = 16'd15;
         684      :	result = 16'd15;
         685      :	result = 16'd15;
         686      :	result = 16'd15;
         687      :	result = 16'd15;
         688      :	result = 16'd15;
         689      :	result = 16'd15;
         690      :	result = 16'd15;
         691      :	result = 16'd15;
         692      :	result = 16'd15;
         693      :	result = 16'd14;
         694      :	result = 16'd14;
         695      :	result = 16'd14;
         696      :	result = 16'd14;
         697      :	result = 16'd14;
         698      :	result = 16'd14;
         699      :	result = 16'd14;
         700      :	result = 16'd14;
         701      :	result = 16'd14;
         702      :	result = 16'd14;
         703      :	result = 16'd14;
         704      :	result = 16'd14;
         705      :	result = 16'd14;
         706      :	result = 16'd14;
         707      :	result = 16'd14;
         708      :	result = 16'd14;
         709      :	result = 16'd14;
         710      :	result = 16'd14;
         711      :	result = 16'd14;
         712      :	result = 16'd14;
         713      :	result = 16'd13;
         714      :	result = 16'd13;
         715      :	result = 16'd13;
         716      :	result = 16'd13;
         717      :	result = 16'd13;
         718      :	result = 16'd13;
         719      :	result = 16'd13;
         720      :	result = 16'd13;
         721      :	result = 16'd13;
         722      :	result = 16'd13;
         723      :	result = 16'd13;
         724      :	result = 16'd13;
         725      :	result = 16'd13;
         726      :	result = 16'd13;
         727      :	result = 16'd13;
         728      :	result = 16'd13;
         729      :	result = 16'd13;
         730      :	result = 16'd13;
         731      :	result = 16'd13;
         732      :	result = 16'd13;
         733      :	result = 16'd13;
         734      :	result = 16'd12;
         735      :	result = 16'd12;
         736      :	result = 16'd12;
         737      :	result = 16'd12;
         738      :	result = 16'd12;
         739      :	result = 16'd12;
         740      :	result = 16'd12;
         741      :	result = 16'd12;
         742      :	result = 16'd12;
         743      :	result = 16'd12;
         744      :	result = 16'd12;
         745      :	result = 16'd12;
         746      :	result = 16'd12;
         747      :	result = 16'd12;
         748      :	result = 16'd12;
         749      :	result = 16'd12;
         750      :	result = 16'd12;
         751      :	result = 16'd12;
         752      :	result = 16'd12;
         753      :	result = 16'd12;
         754      :	result = 16'd12;
         755      :	result = 16'd12;
         756      :	result = 16'd12;
         757      :	result = 16'd11;
         758      :	result = 16'd11;
         759      :	result = 16'd11;
         760      :	result = 16'd11;
         761      :	result = 16'd11;
         762      :	result = 16'd11;
         763      :	result = 16'd11;
         764      :	result = 16'd11;
         765      :	result = 16'd11;
         766      :	result = 16'd11;
         767      :	result = 16'd11;
         768      :	result = 16'd11;
         769      :	result = 16'd11;
         770      :	result = 16'd11;
         771      :	result = 16'd11;
         772      :	result = 16'd11;
         773      :	result = 16'd11;
         774      :	result = 16'd11;
         775      :	result = 16'd11;
         776      :	result = 16'd11;
         777      :	result = 16'd11;
         778      :	result = 16'd11;
         779      :	result = 16'd11;
         780      :	result = 16'd11;
         781      :	result = 16'd11;
         782      :	result = 16'd10;
         783      :	result = 16'd10;
         784      :	result = 16'd10;
         785      :	result = 16'd10;
         786      :	result = 16'd10;
         787      :	result = 16'd10;
         788      :	result = 16'd10;
         789      :	result = 16'd10;
         790      :	result = 16'd10;
         791      :	result = 16'd10;
         792      :	result = 16'd10;
         793      :	result = 16'd10;
         794      :	result = 16'd10;
         795      :	result = 16'd10;
         796      :	result = 16'd10;
         797      :	result = 16'd10;
         798      :	result = 16'd10;
         799      :	result = 16'd10;
         800      :	result = 16'd10;
         801      :	result = 16'd10;
         802      :	result = 16'd10;
         803      :	result = 16'd10;
         804      :	result = 16'd10;
         805      :	result = 16'd10;
         806      :	result = 16'd10;
         807      :	result = 16'd10;
         808      :	result = 16'd9;
         809      :	result = 16'd9;
         810      :	result = 16'd9;
         811      :	result = 16'd9;
         812      :	result = 16'd9;
         813      :	result = 16'd9;
         814      :	result = 16'd9;
         815      :	result = 16'd9;
         816      :	result = 16'd9;
         817      :	result = 16'd9;
         818      :	result = 16'd9;
         819      :	result = 16'd9;
         820      :	result = 16'd9;
         821      :	result = 16'd9;
         822      :	result = 16'd9;
         823      :	result = 16'd9;
         824      :	result = 16'd9;
         825      :	result = 16'd9;
         826      :	result = 16'd9;
         827      :	result = 16'd9;
         828      :	result = 16'd9;
         829      :	result = 16'd9;
         830      :	result = 16'd9;
         831      :	result = 16'd9;
         832      :	result = 16'd9;
         833      :	result = 16'd9;
         834      :	result = 16'd9;
         835      :	result = 16'd9;
         836      :	result = 16'd9;
         837      :	result = 16'd9;
         838      :	result = 16'd8;
         839      :	result = 16'd8;
         840      :	result = 16'd8;
         841      :	result = 16'd8;
         842      :	result = 16'd8;
         843      :	result = 16'd8;
         844      :	result = 16'd8;
         845      :	result = 16'd8;
         846      :	result = 16'd8;
         847      :	result = 16'd8;
         848      :	result = 16'd8;
         849      :	result = 16'd8;
         850      :	result = 16'd8;
         851      :	result = 16'd8;
         852      :	result = 16'd8;
         853      :	result = 16'd8;
         854      :	result = 16'd8;
         855      :	result = 16'd8;
         856      :	result = 16'd8;
         857      :	result = 16'd8;
         858      :	result = 16'd8;
         859      :	result = 16'd8;
         860      :	result = 16'd8;
         861      :	result = 16'd8;
         862      :	result = 16'd8;
         863      :	result = 16'd8;
         864      :	result = 16'd8;
         865      :	result = 16'd8;
         866      :	result = 16'd8;
         867      :	result = 16'd8;
         868      :	result = 16'd8;
         869      :	result = 16'd8;
         870      :	result = 16'd7;
         871      :	result = 16'd7;
         872      :	result = 16'd7;
         873      :	result = 16'd7;
         874      :	result = 16'd7;
         875      :	result = 16'd7;
         876      :	result = 16'd7;
         877      :	result = 16'd7;
         878      :	result = 16'd7;
         879      :	result = 16'd7;
         880      :	result = 16'd7;
         881      :	result = 16'd7;
         882      :	result = 16'd7;
         883      :	result = 16'd7;
         884      :	result = 16'd7;
         885      :	result = 16'd7;
         886      :	result = 16'd7;
         887      :	result = 16'd7;
         888      :	result = 16'd7;
         889      :	result = 16'd7;
         890      :	result = 16'd7;
         891      :	result = 16'd7;
         892      :	result = 16'd7;
         893      :	result = 16'd7;
         894      :	result = 16'd7;
         895      :	result = 16'd7;
         896      :	result = 16'd7;
         897      :	result = 16'd7;
         898      :	result = 16'd7;
         899      :	result = 16'd7;
         900      :	result = 16'd7;
         901      :	result = 16'd7;
         902      :	result = 16'd7;
         903      :	result = 16'd7;
         904      :	result = 16'd7;
         905      :	result = 16'd7;
         906      :	result = 16'd6;
         907      :	result = 16'd6;
         908      :	result = 16'd6;
         909      :	result = 16'd6;
         910      :	result = 16'd6;
         911      :	result = 16'd6;
         912      :	result = 16'd6;
         913      :	result = 16'd6;
         914      :	result = 16'd6;
         915      :	result = 16'd6;
         916      :	result = 16'd6;
         917      :	result = 16'd6;
         918      :	result = 16'd6;
         919      :	result = 16'd6;
         920      :	result = 16'd6;
         921      :	result = 16'd6;
         922      :	result = 16'd6;
         923      :	result = 16'd6;
         924      :	result = 16'd6;
         925      :	result = 16'd6;
         926      :	result = 16'd6;
         927      :	result = 16'd6;
         928      :	result = 16'd6;
         929      :	result = 16'd6;
         930      :	result = 16'd6;
         931      :	result = 16'd6;
         932      :	result = 16'd6;
         933      :	result = 16'd6;
         934      :	result = 16'd6;
         935      :	result = 16'd6;
         936      :	result = 16'd6;
         937      :	result = 16'd6;
         938      :	result = 16'd6;
         939      :	result = 16'd6;
         940      :	result = 16'd6;
         941      :	result = 16'd6;
         942      :	result = 16'd6;
         943      :	result = 16'd6;
         944      :	result = 16'd6;
         945      :	result = 16'd6;
         946      :	result = 16'd6;
         947      :	result = 16'd6;
         948      :	result = 16'd5;
         949      :	result = 16'd5;
         950      :	result = 16'd5;
         951      :	result = 16'd5;
         952      :	result = 16'd5;
         953      :	result = 16'd5;
         954      :	result = 16'd5;
         955      :	result = 16'd5;
         956      :	result = 16'd5;
         957      :	result = 16'd5;
         958      :	result = 16'd5;
         959      :	result = 16'd5;
         960      :	result = 16'd5;
         961      :	result = 16'd5;
         962      :	result = 16'd5;
         963      :	result = 16'd5;
         964      :	result = 16'd5;
         965      :	result = 16'd5;
         966      :	result = 16'd5;
         967      :	result = 16'd5;
         968      :	result = 16'd5;
         969      :	result = 16'd5;
         970      :	result = 16'd5;
         971      :	result = 16'd5;
         972      :	result = 16'd5;
         973      :	result = 16'd5;
         974      :	result = 16'd5;
         975      :	result = 16'd5;
         976      :	result = 16'd5;
         977      :	result = 16'd5;
         978      :	result = 16'd5;
         979      :	result = 16'd5;
         980      :	result = 16'd5;
         981      :	result = 16'd5;
         982      :	result = 16'd5;
         983      :	result = 16'd5;
         984      :	result = 16'd5;
         985      :	result = 16'd5;
         986      :	result = 16'd5;
         987      :	result = 16'd5;
         988      :	result = 16'd5;
         989      :	result = 16'd5;
         990      :	result = 16'd5;
         991      :	result = 16'd5;
         992      :	result = 16'd5;
         993      :	result = 16'd5;
         994      :	result = 16'd5;
         995      :	result = 16'd5;
         996      :	result = 16'd5;
         997      :	result = 16'd4;
         998      :	result = 16'd4;
         999      :	result = 16'd4;
         1000     :	result = 16'd4;
         1001     :	result = 16'd4;
         1002     :	result = 16'd4;
         1003     :	result = 16'd4;
         1004     :	result = 16'd4;
         1005     :	result = 16'd4;
         1006     :	result = 16'd4;
         1007     :	result = 16'd4;
         1008     :	result = 16'd4;
         1009     :	result = 16'd4;
         1010     :	result = 16'd4;
         1011     :	result = 16'd4;
         1012     :	result = 16'd4;
         1013     :	result = 16'd4;
         1014     :	result = 16'd4;
         1015     :	result = 16'd4;
         1016     :	result = 16'd4;
         1017     :	result = 16'd4;
         1018     :	result = 16'd4;
         1019     :	result = 16'd4;
         1020     :	result = 16'd4;
         1021     :	result = 16'd4;
         1022     :	result = 16'd4;
         1023     :	result = 16'd4;
         1024     :	result = 16'd4;
         1025     :	result = 16'd4;
         1026     :	result = 16'd4;
         1027     :	result = 16'd4;
         1028     :	result = 16'd4;
         1029     :	result = 16'd4;
         1030     :	result = 16'd4;
         1031     :	result = 16'd4;
         1032     :	result = 16'd4;
         1033     :	result = 16'd4;
         1034     :	result = 16'd4;
         1035     :	result = 16'd4;
         1036     :	result = 16'd4;
         1037     :	result = 16'd4;
         1038     :	result = 16'd4;
         1039     :	result = 16'd4;
         1040     :	result = 16'd4;
         1041     :	result = 16'd4;
         1042     :	result = 16'd4;
         1043     :	result = 16'd4;
         1044     :	result = 16'd4;
         1045     :	result = 16'd4;
         1046     :	result = 16'd4;
         1047     :	result = 16'd4;
         1048     :	result = 16'd4;
         1049     :	result = 16'd4;
         1050     :	result = 16'd4;
         1051     :	result = 16'd4;
         1052     :	result = 16'd4;
         1053     :	result = 16'd4;
         1054     :	result = 16'd4;
         1055     :	result = 16'd4;
         1056     :	result = 16'd3;
         1057     :	result = 16'd3;
         1058     :	result = 16'd3;
         1059     :	result = 16'd3;
         1060     :	result = 16'd3;
         1061     :	result = 16'd3;
         1062     :	result = 16'd3;
         1063     :	result = 16'd3;
         1064     :	result = 16'd3;
         1065     :	result = 16'd3;
         1066     :	result = 16'd3;
         1067     :	result = 16'd3;
         1068     :	result = 16'd3;
         1069     :	result = 16'd3;
         1070     :	result = 16'd3;
         1071     :	result = 16'd3;
         1072     :	result = 16'd3;
         1073     :	result = 16'd3;
         1074     :	result = 16'd3;
         1075     :	result = 16'd3;
         1076     :	result = 16'd3;
         1077     :	result = 16'd3;
         1078     :	result = 16'd3;
         1079     :	result = 16'd3;
         1080     :	result = 16'd3;
         1081     :	result = 16'd3;
         1082     :	result = 16'd3;
         1083     :	result = 16'd3;
         1084     :	result = 16'd3;
         1085     :	result = 16'd3;
         1086     :	result = 16'd3;
         1087     :	result = 16'd3;
         1088     :	result = 16'd3;
         1089     :	result = 16'd3;
         1090     :	result = 16'd3;
         1091     :	result = 16'd3;
         1092     :	result = 16'd3;
         1093     :	result = 16'd3;
         1094     :	result = 16'd3;
         1095     :	result = 16'd3;
         1096     :	result = 16'd3;
         1097     :	result = 16'd3;
         1098     :	result = 16'd3;
         1099     :	result = 16'd3;
         1100     :	result = 16'd3;
         1101     :	result = 16'd3;
         1102     :	result = 16'd3;
         1103     :	result = 16'd3;
         1104     :	result = 16'd3;
         1105     :	result = 16'd3;
         1106     :	result = 16'd3;
         1107     :	result = 16'd3;
         1108     :	result = 16'd3;
         1109     :	result = 16'd3;
         1110     :	result = 16'd3;
         1111     :	result = 16'd3;
         1112     :	result = 16'd3;
         1113     :	result = 16'd3;
         1114     :	result = 16'd3;
         1115     :	result = 16'd3;
         1116     :	result = 16'd3;
         1117     :	result = 16'd3;
         1118     :	result = 16'd3;
         1119     :	result = 16'd3;
         1120     :	result = 16'd3;
         1121     :	result = 16'd3;
         1122     :	result = 16'd3;
         1123     :	result = 16'd3;
         1124     :	result = 16'd3;
         1125     :	result = 16'd3;
         1126     :	result = 16'd3;
         1127     :	result = 16'd3;
         1128     :	result = 16'd3;
         1129     :	result = 16'd3;
         1130     :	result = 16'd3;
         1131     :	result = 16'd3;
         1132     :	result = 16'd2;
         1133     :	result = 16'd2;
         1134     :	result = 16'd2;
         1135     :	result = 16'd2;
         1136     :	result = 16'd2;
         1137     :	result = 16'd2;
         1138     :	result = 16'd2;
         1139     :	result = 16'd2;
         1140     :	result = 16'd2;
         1141     :	result = 16'd2;
         1142     :	result = 16'd2;
         1143     :	result = 16'd2;
         1144     :	result = 16'd2;
         1145     :	result = 16'd2;
         1146     :	result = 16'd2;
         1147     :	result = 16'd2;
         1148     :	result = 16'd2;
         1149     :	result = 16'd2;
         1150     :	result = 16'd2;
         1151     :	result = 16'd2;
         1152     :	result = 16'd2;
         1153     :	result = 16'd2;
         1154     :	result = 16'd2;
         1155     :	result = 16'd2;
         1156     :	result = 16'd2;
         1157     :	result = 16'd2;
         1158     :	result = 16'd2;
         1159     :	result = 16'd2;
         1160     :	result = 16'd2;
         1161     :	result = 16'd2;
         1162     :	result = 16'd2;
         1163     :	result = 16'd2;
         1164     :	result = 16'd2;
         1165     :	result = 16'd2;
         1166     :	result = 16'd2;
         1167     :	result = 16'd2;
         1168     :	result = 16'd2;
         1169     :	result = 16'd2;
         1170     :	result = 16'd2;
         1171     :	result = 16'd2;
         1172     :	result = 16'd2;
         1173     :	result = 16'd2;
         1174     :	result = 16'd2;
         1175     :	result = 16'd2;
         1176     :	result = 16'd2;
         1177     :	result = 16'd2;
         1178     :	result = 16'd2;
         1179     :	result = 16'd2;
         1180     :	result = 16'd2;
         1181     :	result = 16'd2;
         1182     :	result = 16'd2;
         1183     :	result = 16'd2;
         1184     :	result = 16'd2;
         1185     :	result = 16'd2;
         1186     :	result = 16'd2;
         1187     :	result = 16'd2;
         1188     :	result = 16'd2;
         1189     :	result = 16'd2;
         1190     :	result = 16'd2;
         1191     :	result = 16'd2;
         1192     :	result = 16'd2;
         1193     :	result = 16'd2;
         1194     :	result = 16'd2;
         1195     :	result = 16'd2;
         1196     :	result = 16'd2;
         1197     :	result = 16'd2;
         1198     :	result = 16'd2;
         1199     :	result = 16'd2;
         1200     :	result = 16'd2;
         1201     :	result = 16'd2;
         1202     :	result = 16'd2;
         1203     :	result = 16'd2;
         1204     :	result = 16'd2;
         1205     :	result = 16'd2;
         1206     :	result = 16'd2;
         1207     :	result = 16'd2;
         1208     :	result = 16'd2;
         1209     :	result = 16'd2;
         1210     :	result = 16'd2;
         1211     :	result = 16'd2;
         1212     :	result = 16'd2;
         1213     :	result = 16'd2;
         1214     :	result = 16'd2;
         1215     :	result = 16'd2;
         1216     :	result = 16'd2;
         1217     :	result = 16'd2;
         1218     :	result = 16'd2;
         1219     :	result = 16'd2;
         1220     :	result = 16'd2;
         1221     :	result = 16'd2;
         1222     :	result = 16'd2;
         1223     :	result = 16'd2;
         1224     :	result = 16'd2;
         1225     :	result = 16'd2;
         1226     :	result = 16'd2;
         1227     :	result = 16'd2;
         1228     :	result = 16'd2;
         1229     :	result = 16'd2;
         1230     :	result = 16'd2;
         1231     :	result = 16'd2;
         1232     :	result = 16'd2;
         1233     :	result = 16'd2;
         1234     :	result = 16'd2;
         1235     :	result = 16'd2;
         1236     :	result = 16'd2;
         1237     :	result = 16'd2;
         1238     :	result = 16'd1;
         1239     :	result = 16'd1;
         1240     :	result = 16'd1;
         1241     :	result = 16'd1;
         1242     :	result = 16'd1;
         1243     :	result = 16'd1;
         1244     :	result = 16'd1;
         1245     :	result = 16'd1;
         1246     :	result = 16'd1;
         1247     :	result = 16'd1;
         1248     :	result = 16'd1;
         1249     :	result = 16'd1;
         1250     :	result = 16'd1;
         1251     :	result = 16'd1;
         1252     :	result = 16'd1;
         1253     :	result = 16'd1;
         1254     :	result = 16'd1;
         1255     :	result = 16'd1;
         1256     :	result = 16'd1;
         1257     :	result = 16'd1;
         1258     :	result = 16'd1;
         1259     :	result = 16'd1;
         1260     :	result = 16'd1;
         1261     :	result = 16'd1;
         1262     :	result = 16'd1;
         1263     :	result = 16'd1;
         1264     :	result = 16'd1;
         1265     :	result = 16'd1;
         1266     :	result = 16'd1;
         1267     :	result = 16'd1;
         1268     :	result = 16'd1;
         1269     :	result = 16'd1;
         1270     :	result = 16'd1;
         1271     :	result = 16'd1;
         1272     :	result = 16'd1;
         1273     :	result = 16'd1;
         1274     :	result = 16'd1;
         1275     :	result = 16'd1;
         1276     :	result = 16'd1;
         1277     :	result = 16'd1;
         1278     :	result = 16'd1;
         1279     :	result = 16'd1;
         1280     :	result = 16'd1;
         1281     :	result = 16'd1;
         1282     :	result = 16'd1;
         1283     :	result = 16'd1;
         1284     :	result = 16'd1;
         1285     :	result = 16'd1;
         1286     :	result = 16'd1;
         1287     :	result = 16'd1;
         1288     :	result = 16'd1;
         1289     :	result = 16'd1;
         1290     :	result = 16'd1;
         1291     :	result = 16'd1;
         1292     :	result = 16'd1;
         1293     :	result = 16'd1;
         1294     :	result = 16'd1;
         1295     :	result = 16'd1;
         1296     :	result = 16'd1;
         1297     :	result = 16'd1;
         1298     :	result = 16'd1;
         1299     :	result = 16'd1;
         1300     :	result = 16'd1;
         1301     :	result = 16'd1;
         1302     :	result = 16'd1;
         1303     :	result = 16'd1;
         1304     :	result = 16'd1;
         1305     :	result = 16'd1;
         1306     :	result = 16'd1;
         1307     :	result = 16'd1;
         1308     :	result = 16'd1;
         1309     :	result = 16'd1;
         1310     :	result = 16'd1;
         1311     :	result = 16'd1;
         1312     :	result = 16'd1;
         1313     :	result = 16'd1;
         1314     :	result = 16'd1;
         1315     :	result = 16'd1;
         1316     :	result = 16'd1;
         1317     :	result = 16'd1;
         1318     :	result = 16'd1;
         1319     :	result = 16'd1;
         1320     :	result = 16'd1;
         1321     :	result = 16'd1;
         1322     :	result = 16'd1;
         1323     :	result = 16'd1;
         1324     :	result = 16'd1;
         1325     :	result = 16'd1;
         1326     :	result = 16'd1;
         1327     :	result = 16'd1;
         1328     :	result = 16'd1;
         1329     :	result = 16'd1;
         1330     :	result = 16'd1;
         1331     :	result = 16'd1;
         1332     :	result = 16'd1;
         1333     :	result = 16'd1;
         1334     :	result = 16'd1;
         1335     :	result = 16'd1;
         1336     :	result = 16'd1;
         1337     :	result = 16'd1;
         1338     :	result = 16'd1;
         1339     :	result = 16'd1;
         1340     :	result = 16'd1;
         1341     :	result = 16'd1;
         1342     :	result = 16'd1;
         1343     :	result = 16'd1;
         1344     :	result = 16'd1;
         1345     :	result = 16'd1;
         1346     :	result = 16'd1;
         1347     :	result = 16'd1;
         1348     :	result = 16'd1;
         1349     :	result = 16'd1;
         1350     :	result = 16'd1;
         1351     :	result = 16'd1;
         1352     :	result = 16'd1;
         1353     :	result = 16'd1;
         1354     :	result = 16'd1;
         1355     :	result = 16'd1;
         1356     :	result = 16'd1;
         1357     :	result = 16'd1;
         1358     :	result = 16'd1;
         1359     :	result = 16'd1;
         1360     :	result = 16'd1;
         1361     :	result = 16'd1;
         1362     :	result = 16'd1;
         1363     :	result = 16'd1;
         1364     :	result = 16'd1;
         1365     :	result = 16'd1;
         1366     :	result = 16'd1;
         1367     :	result = 16'd1;
         1368     :	result = 16'd1;
         1369     :	result = 16'd1;
         1370     :	result = 16'd1;
         1371     :	result = 16'd1;
         1372     :	result = 16'd1;
         1373     :	result = 16'd1;
         1374     :	result = 16'd1;
         1375     :	result = 16'd1;
         1376     :	result = 16'd1;
         1377     :	result = 16'd1;
         1378     :	result = 16'd1;
         1379     :	result = 16'd1;
         1380     :	result = 16'd1;
         1381     :	result = 16'd1;
         1382     :	result = 16'd1;
         1383     :	result = 16'd1;
         1384     :	result = 16'd1;
         1385     :	result = 16'd1;
         1386     :	result = 16'd1;
         1387     :	result = 16'd1;
         1388     :	result = 16'd1;
         1389     :	result = 16'd1;
         1390     :	result = 16'd1;
         1391     :	result = 16'd1;
         1392     :	result = 16'd1;
         1393     :	result = 16'd1;
         1394     :	result = 16'd1;
         1395     :	result = 16'd1;
         1396     :	result = 16'd1;
         1397     :	result = 16'd1;
         1398     :	result = 16'd1;
         1399     :	result = 16'd1;
         1400     :	result = 16'd1;
         1401     :	result = 16'd1;
         1402     :	result = 16'd1;
         1403     :	result = 16'd1;
         1404     :	result = 16'd1;
         1405     :	result = 16'd1;
         1406     :	result = 16'd1;
         1407     :	result = 16'd1;
         1408     :	result = 16'd1;
         1409     :	result = 16'd1;
         1410     :	result = 16'd1;
         1411     :	result = 16'd1;
         1412     :	result = 16'd1;
         1413     :	result = 16'd1;
         1414     :	result = 16'd1;
         1415     :	result = 16'd1;
         1416     :	result = 16'd1;
         1417     :	result = 16'd0;
         1418     :	result = 16'd0;
         1419     :	result = 16'd0;
         1420     :	result = 16'd0;
         1421     :	result = 16'd0;
         1422     :	result = 16'd0;
         1423     :	result = 16'd0;
         1424     :	result = 16'd0;
         1425     :	result = 16'd0;
         1426     :	result = 16'd0;
         1427     :	result = 16'd0;
         1428     :	result = 16'd0;
         1429     :	result = 16'd0;
         1430     :	result = 16'd0;
         1431     :	result = 16'd0;
         1432     :	result = 16'd0;
         1433     :	result = 16'd0;
         1434     :	result = 16'd0;
         1435     :	result = 16'd0;
         1436     :	result = 16'd0;
         1437     :	result = 16'd0;
         1438     :	result = 16'd0;
         1439     :	result = 16'd0;
         1440     :	result = 16'd0;
         1441     :	result = 16'd0;
         1442     :	result = 16'd0;
         1443     :	result = 16'd0;
         1444     :	result = 16'd0;
         1445     :	result = 16'd0;
         1446     :	result = 16'd0;
         1447     :	result = 16'd0;
         1448     :	result = 16'd0;
         1449     :	result = 16'd0;
         1450     :	result = 16'd0;
         1451     :	result = 16'd0;
         1452     :	result = 16'd0;
         1453     :	result = 16'd0;
         1454     :	result = 16'd0;
         1455     :	result = 16'd0;
         1456     :	result = 16'd0;
         1457     :	result = 16'd0;
         1458     :	result = 16'd0;
         1459     :	result = 16'd0;
         1460     :	result = 16'd0;
         1461     :	result = 16'd0;
         1462     :	result = 16'd0;
         1463     :	result = 16'd0;
         1464     :	result = 16'd0;
         1465     :	result = 16'd0;
         1466     :	result = 16'd0;
         1467     :	result = 16'd0;
         1468     :	result = 16'd0;
         1469     :	result = 16'd0;
         1470     :	result = 16'd0;
         1471     :	result = 16'd0;
         1472     :	result = 16'd0;
         1473     :	result = 16'd0;
         1474     :	result = 16'd0;
         1475     :	result = 16'd0;
         1476     :	result = 16'd0;
         1477     :	result = 16'd0;
         1478     :	result = 16'd0;
         1479     :	result = 16'd0;
         1480     :	result = 16'd0;
         1481     :	result = 16'd0;
         1482     :	result = 16'd0;
         1483     :	result = 16'd0;
         1484     :	result = 16'd0;
         1485     :	result = 16'd0;
         1486     :	result = 16'd0;
         1487     :	result = 16'd0;
         1488     :	result = 16'd0;
         1489     :	result = 16'd0;
         1490     :	result = 16'd0;
         1491     :	result = 16'd0;
         1492     :	result = 16'd0;
         1493     :	result = 16'd0;
         1494     :	result = 16'd0;
         1495     :	result = 16'd0;
         1496     :	result = 16'd0;
         1497     :	result = 16'd0;
         1498     :	result = 16'd0;
         1499     :	result = 16'd0;
         1500     :	result = 16'd0;
         1501     :	result = 16'd0;
         1502     :	result = 16'd0;
         1503     :	result = 16'd0;
         1504     :	result = 16'd0;
         1505     :	result = 16'd0;
         1506     :	result = 16'd0;
         1507     :	result = 16'd0;
         1508     :	result = 16'd0;
         1509     :	result = 16'd0;
         1510     :	result = 16'd0;
         1511     :	result = 16'd0;
         1512     :	result = 16'd0;
         1513     :	result = 16'd0;
         1514     :	result = 16'd0;
         1515     :	result = 16'd0;
         1516     :	result = 16'd0;
         1517     :	result = 16'd0;
         1518     :	result = 16'd0;
         1519     :	result = 16'd0;
         1520     :	result = 16'd0;
         1521     :	result = 16'd0;
         1522     :	result = 16'd0;
         1523     :	result = 16'd0;
         1524     :	result = 16'd0;
         1525     :	result = 16'd0;
         1526     :	result = 16'd0;
         1527     :	result = 16'd0;
         1528     :	result = 16'd0;
         1529     :	result = 16'd0;
         1530     :	result = 16'd0;
         1531     :	result = 16'd0;
         1532     :	result = 16'd0;
         1533     :	result = 16'd0;
         1534     :	result = 16'd0;
         1535     :	result = 16'd0;
         1536     :	result = 16'd0;
         1537     :	result = 16'd0;
         1538     :	result = 16'd0;
         1539     :	result = 16'd0;
         1540     :	result = 16'd0;
         1541     :	result = 16'd0;
         1542     :	result = 16'd0;
         1543     :	result = 16'd0;
         1544     :	result = 16'd0;
         1545     :	result = 16'd0;
         1546     :	result = 16'd0;
         1547     :	result = 16'd0;
         1548     :	result = 16'd0;
         1549     :	result = 16'd0;
         1550     :	result = 16'd0;
         1551     :	result = 16'd0;
         1552     :	result = 16'd0;
         1553     :	result = 16'd0;
         1554     :	result = 16'd0;
         1555     :	result = 16'd0;
         1556     :	result = 16'd0;
         1557     :	result = 16'd0;
         1558     :	result = 16'd0;
         1559     :	result = 16'd0;
         1560     :	result = 16'd0;
         1561     :	result = 16'd0;
         1562     :	result = 16'd0;
         1563     :	result = 16'd0;
         1564     :	result = 16'd0;
         1565     :	result = 16'd0;
         1566     :	result = 16'd0;
         1567     :	result = 16'd0;
         1568     :	result = 16'd0;
         1569     :	result = 16'd0;
         1570     :	result = 16'd0;
         1571     :	result = 16'd0;
         1572     :	result = 16'd0;
         1573     :	result = 16'd0;
         1574     :	result = 16'd0;
         1575     :	result = 16'd0;
         1576     :	result = 16'd0;
         1577     :	result = 16'd0;
         1578     :	result = 16'd0;
         1579     :	result = 16'd0;
         1580     :	result = 16'd0;
         1581     :	result = 16'd0;
         1582     :	result = 16'd0;
         1583     :	result = 16'd0;
         1584     :	result = 16'd0;
         1585     :	result = 16'd0;
         1586     :	result = 16'd0;
         1587     :	result = 16'd0;
         1588     :	result = 16'd0;
         1589     :	result = 16'd0;
         1590     :	result = 16'd0;
         1591     :	result = 16'd0;
         1592     :	result = 16'd0;
         1593     :	result = 16'd0;
         1594     :	result = 16'd0;
         1595     :	result = 16'd0;
         1596     :	result = 16'd0;
         1597     :	result = 16'd0;
         1598     :	result = 16'd0;
         1599     :	result = 16'd0;
         1600     :	result = 16'd0;
         1601     :	result = 16'd0;
         1602     :	result = 16'd0;
         1603     :	result = 16'd0;
         1604     :	result = 16'd0;
         1605     :	result = 16'd0;
         1606     :	result = 16'd0;
         1607     :	result = 16'd0;
         1608     :	result = 16'd0;
         1609     :	result = 16'd0;
         1610     :	result = 16'd0;
         1611     :	result = 16'd0;
         1612     :	result = 16'd0;
         1613     :	result = 16'd0;
         1614     :	result = 16'd0;
         1615     :	result = 16'd0;
         1616     :	result = 16'd0;
         1617     :	result = 16'd0;
         1618     :	result = 16'd0;
         1619     :	result = 16'd0;
         1620     :	result = 16'd0;
         1621     :	result = 16'd0;
         1622     :	result = 16'd0;
         1623     :	result = 16'd0;
         1624     :	result = 16'd0;
         1625     :	result = 16'd0;
         1626     :	result = 16'd0;
         1627     :	result = 16'd0;
         1628     :	result = 16'd0;
         1629     :	result = 16'd0;
         1630     :	result = 16'd0;
         1631     :	result = 16'd0;
         1632     :	result = 16'd0;
         1633     :	result = 16'd0;
         1634     :	result = 16'd0;
         1635     :	result = 16'd0;
         1636     :	result = 16'd0;
         1637     :	result = 16'd0;
         1638     :	result = 16'd0;
         1639     :	result = 16'd0;
         1640     :	result = 16'd0;
         1641     :	result = 16'd0;
         1642     :	result = 16'd0;
         1643     :	result = 16'd0;
         1644     :	result = 16'd0;
         1645     :	result = 16'd0;
         1646     :	result = 16'd0;
         1647     :	result = 16'd0;
         1648     :	result = 16'd0;
         1649     :	result = 16'd0;
         1650     :	result = 16'd0;
         1651     :	result = 16'd0;
         1652     :	result = 16'd0;
         1653     :	result = 16'd0;
         1654     :	result = 16'd0;
         1655     :	result = 16'd0;
         1656     :	result = 16'd0;
         1657     :	result = 16'd0;
         1658     :	result = 16'd0;
         1659     :	result = 16'd0;
         1660     :	result = 16'd0;
         1661     :	result = 16'd0;
         1662     :	result = 16'd0;
         1663     :	result = 16'd0;
         1664     :	result = 16'd0;
         1665     :	result = 16'd0;
         1666     :	result = 16'd0;
         1667     :	result = 16'd0;
         1668     :	result = 16'd0;
         1669     :	result = 16'd0;
         1670     :	result = 16'd0;
         1671     :	result = 16'd0;
         1672     :	result = 16'd0;
         1673     :	result = 16'd0;
         1674     :	result = 16'd0;
         1675     :	result = 16'd0;
         1676     :	result = 16'd0;
         1677     :	result = 16'd0;
         1678     :	result = 16'd0;
         1679     :	result = 16'd0;
         1680     :	result = 16'd0;
         1681     :	result = 16'd0;
         1682     :	result = 16'd0;
         1683     :	result = 16'd0;
         1684     :	result = 16'd0;
         1685     :	result = 16'd0;
         1686     :	result = 16'd0;
         1687     :	result = 16'd0;
         1688     :	result = 16'd0;
         1689     :	result = 16'd0;
         1690     :	result = 16'd0;
         1691     :	result = 16'd0;
         1692     :	result = 16'd0;
         1693     :	result = 16'd0;
         1694     :	result = 16'd0;
         1695     :	result = 16'd0;
         1696     :	result = 16'd0;
         1697     :	result = 16'd0;
         1698     :	result = 16'd0;
         1699     :	result = 16'd0;
         1700     :	result = 16'd0;
         1701     :	result = 16'd0;
         1702     :	result = 16'd0;
         1703     :	result = 16'd0;
         1704     :	result = 16'd0;
         1705     :	result = 16'd0;
         1706     :	result = 16'd0;
         1707     :	result = 16'd0;
         1708     :	result = 16'd0;
         1709     :	result = 16'd0;
         1710     :	result = 16'd0;
         1711     :	result = 16'd0;
         1712     :	result = 16'd0;
         1713     :	result = 16'd0;
         1714     :	result = 16'd0;
         1715     :	result = 16'd0;
         1716     :	result = 16'd0;
         1717     :	result = 16'd0;
         1718     :	result = 16'd0;
         1719     :	result = 16'd0;
         1720     :	result = 16'd0;
         1721     :	result = 16'd0;
         1722     :	result = 16'd0;
         1723     :	result = 16'd0;
         1724     :	result = 16'd0;
         1725     :	result = 16'd0;
         1726     :	result = 16'd0;
         1727     :	result = 16'd0;
         1728     :	result = 16'd0;
         1729     :	result = 16'd0;
         1730     :	result = 16'd0;
         1731     :	result = 16'd0;
         1732     :	result = 16'd0;
         1733     :	result = 16'd0;
         1734     :	result = 16'd0;
         1735     :	result = 16'd0;
         1736     :	result = 16'd0;
         1737     :	result = 16'd0;
         1738     :	result = 16'd0;
         1739     :	result = 16'd0;
         1740     :	result = 16'd0;
         1741     :	result = 16'd0;
         1742     :	result = 16'd0;
         1743     :	result = 16'd0;
         1744     :	result = 16'd0;
         1745     :	result = 16'd0;
         1746     :	result = 16'd0;
         1747     :	result = 16'd0;
         1748     :	result = 16'd0;
         1749     :	result = 16'd0;
         1750     :	result = 16'd0;
         1751     :	result = 16'd0;
         1752     :	result = 16'd0;
         1753     :	result = 16'd0;
         1754     :	result = 16'd0;
         1755     :	result = 16'd0;
         1756     :	result = 16'd0;
         1757     :	result = 16'd0;
         1758     :	result = 16'd0;
         1759     :	result = 16'd0;
         1760     :	result = 16'd0;
         1761     :	result = 16'd0;
         1762     :	result = 16'd0;
         1763     :	result = 16'd0;
         1764     :	result = 16'd0;
         1765     :	result = 16'd0;
         1766     :	result = 16'd0;
         1767     :	result = 16'd0;
         1768     :	result = 16'd0;
         1769     :	result = 16'd0;
         1770     :	result = 16'd0;
         1771     :	result = 16'd0;
         1772     :	result = 16'd0;
         1773     :	result = 16'd0;
         1774     :	result = 16'd0;
         1775     :	result = 16'd0;
         1776     :	result = 16'd0;
         1777     :	result = 16'd0;
         1778     :	result = 16'd0;
         1779     :	result = 16'd0;
         1780     :	result = 16'd0;
         1781     :	result = 16'd0;
         1782     :	result = 16'd0;
         1783     :	result = 16'd0;
         1784     :	result = 16'd0;
         1785     :	result = 16'd0;
         1786     :	result = 16'd0;
         1787     :	result = 16'd0;
         1788     :	result = 16'd0;
         1789     :	result = 16'd0;
         1790     :	result = 16'd0;
         1791     :	result = 16'd0;
         default  :  result = 16'd0;
      endcase
   end

endmodule